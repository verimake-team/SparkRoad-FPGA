// Verilog netlist created by TD v4.3.815
// Tue May 14 16:19:40 2019

`timescale 1ns / 1ps
module system  // ../src/top.v(3)
  (
  clk,
  resetn_i,
  rxd,
  out_byte,
  out_byte_en,
  trap,
  txd
  );

  input clk;  // ../src/top.v(4)
  input resetn_i;  // ../src/top.v(5)
  input rxd;  // ../src/top.v(14)
  output [7:0] out_byte;  // ../src/top.v(7)
  output out_byte_en;  // ../src/top.v(8)
  output trap;  // ../src/top.v(6)
  output txd;  // ../src/top.v(13)

  wire [1:0] initial_reset;  // ../src/top.v(34)
  wire [31:0] mem_la_addr;  // ../src/top.v(29)
  wire [31:0] mem_la_wdata;  // ../src/top.v(30)
  wire [31:0] mem_rdata;  // ../src/top.v(23)
  wire [31:0] memory_out;  // ../src/top.v(66)
  wire [7:0] n17;
  wire [31:0] \picorv32_core/alu_out_q ;  // ../src/picorv32.v(1174)
  wire [63:0] \picorv32_core/count_cycle ;  // ../src/picorv32.v(145)
  wire [63:0] \picorv32_core/count_instr ;  // ../src/picorv32.v(145)
  wire [7:0] \picorv32_core/cpu_state ;  // ../src/picorv32.v(1134)
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c0_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c0_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c1_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c1_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c2_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c2_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c3_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c3_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c4_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c4_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c5_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c5_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c6_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c6_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c7_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r0_c7_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c0_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c0_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c1_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c1_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c2_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c2_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c3_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c3_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c4_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c4_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c5_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c5_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c6_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c6_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c7_di ;
  wire [3:0] \picorv32_core/cpuregs_p1/dram_r1_c7_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c0_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c0_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c1_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c1_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c2_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c2_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c3_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c3_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c4_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c4_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c5_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c5_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c6_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c6_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c7_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r0_c7_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c0_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c0_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c1_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c1_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c2_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c2_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c3_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c3_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c4_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c4_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c5_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c5_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c6_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c6_waddr ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c7_di ;
  wire [3:0] \picorv32_core/cpuregs_p2/dram_r1_c7_waddr ;
  wire [31:0] \picorv32_core/cpuregs_rs2 ;  // ../src/picorv32.v(1255)
  wire [31:0] \picorv32_core/cpuregs_wrdata ;  // ../src/picorv32.v(1252)
  wire [31:0] \picorv32_core/decoded_imm ;  // ../src/picorv32.v(620)
  wire [31:0] \picorv32_core/decoded_imm_uj ;  // ../src/picorv32.v(620)
  wire [4:0] \picorv32_core/decoded_rd ;  // ../src/picorv32.v(619)
  wire [4:0] \picorv32_core/decoded_rs1 ;  // ../src/picorv32.v(619)
  wire [4:0] \picorv32_core/decoded_rs2 ;  // ../src/picorv32.v(619)
  wire [4:0] \picorv32_core/latched_rd ;  // ../src/picorv32.v(1163)
  wire [15:0] \picorv32_core/mem_16bit_buffer ;  // ../src/picorv32.v(331)
  wire [31:0] \picorv32_core/mem_rdata_latched ;  // ../src/picorv32.v(334)
  wire [31:0] \picorv32_core/mem_rdata_latched_noshuffle ;  // ../src/picorv32.v(333)
  wire [31:0] \picorv32_core/mem_rdata_q ;  // ../src/picorv32.v(319)
  wire [1:0] \picorv32_core/mem_state ;  // ../src/picorv32.v(316)
  wire [1:0] \picorv32_core/mem_wordsize ;  // ../src/picorv32.v(317)
  wire  \picorv32_core/mux79_b0/B0_3 ;
  wire  \picorv32_core/mux79_b0/B1_0 ;
  wire  \picorv32_core/mux79_b1/B0_3 ;
  wire  \picorv32_core/mux79_b2/B0_3 ;
  wire  \picorv32_core/mux79_b3/B1_0 ;
  wire [29:0] \picorv32_core/n30 ;
  wire [3:0] \picorv32_core/n40 ;
  wire [31:0] \picorv32_core/n42 ;
  wire [31:0] \picorv32_core/n433 ;
  wire [31:0] \picorv32_core/n434 ;
  wire [2:0] \picorv32_core/n449 ;
  wire [31:0] \picorv32_core/n450 ;
  wire [63:0] \picorv32_core/n459 ;
  wire [31:0] \picorv32_core/n500 ;
  wire [2:0] \picorv32_core/n501 ;
  wire [31:0] \picorv32_core/n502 ;
  wire [63:0] \picorv32_core/n503 ;
  wire [31:0] \picorv32_core/n504 ;
  wire [7:0] \picorv32_core/n524 ;
  wire [31:0] \picorv32_core/n543 ;
  wire [5:0] \picorv32_core/n559 ;
  wire [5:0] \picorv32_core/n564 ;
  wire [31:0] \picorv32_core/n570 ;
  wire [31:0] \picorv32_core/n576 ;
  wire [2:0] \picorv32_core/n68 ;
  wire [31:0] \picorv32_core/next_pc ;  // ../src/picorv32.v(168)
  wire [31:0] \picorv32_core/reg_next_pc ;  // ../src/picorv32.v(146)
  wire [31:0] \picorv32_core/reg_out ;  // ../src/picorv32.v(146)
  wire [31:0] \picorv32_core/reg_pc ;  // ../src/picorv32.v(146)
  wire [4:0] \picorv32_core/reg_sh ;  // ../src/picorv32.v(151)
  wire  \picorv32_core/sel10_b0/B1_1 ;
  wire  \picorv32_core/sel10_b1/B1_1 ;
  wire  \picorv32_core/sel10_b2/B1_1 ;
  wire  \picorv32_core/sel10_b3/B1_1 ;
  wire  \picorv32_core/sel23/B2 ;
  wire  \picorv32_core/sel27_b16/B1 ;
  wire  \picorv32_core/sel27_b16/B2 ;
  wire  \picorv32_core/sel27_b17/B2 ;
  wire  \picorv32_core/sel27_b18/B2 ;
  wire  \picorv32_core/sel27_b19/B2 ;
  wire  \picorv32_core/sel27_b20/B2 ;
  wire  \picorv32_core/sel27_b21/B2 ;
  wire  \picorv32_core/sel27_b22/B2 ;
  wire  \picorv32_core/sel27_b23/B2 ;
  wire  \picorv32_core/sel27_b24/B2 ;
  wire  \picorv32_core/sel27_b25/B2 ;
  wire  \picorv32_core/sel27_b26/B2 ;
  wire  \picorv32_core/sel27_b27/B2 ;
  wire  \picorv32_core/sel27_b28/B2 ;
  wire  \picorv32_core/sel27_b29/B2 ;
  wire  \picorv32_core/sel27_b30/B2 ;
  wire  \picorv32_core/sel27_b31/B2 ;
  wire  \picorv32_core/sel40_b6/B3 ;
  wire  \picorv32_core/sel40_b6/B5 ;
  wire  \picorv32_core/sel41_b0/B5 ;
  wire  \picorv32_core/sel41_b1/B5 ;
  wire  \picorv32_core/sel41_b10/B2 ;
  wire  \picorv32_core/sel41_b10/B5 ;
  wire  \picorv32_core/sel41_b11/B2 ;
  wire  \picorv32_core/sel41_b11/B5 ;
  wire  \picorv32_core/sel41_b12/B2 ;
  wire  \picorv32_core/sel41_b12/B5 ;
  wire  \picorv32_core/sel41_b13/B2 ;
  wire  \picorv32_core/sel41_b13/B5 ;
  wire  \picorv32_core/sel41_b14/B2 ;
  wire  \picorv32_core/sel41_b14/B5 ;
  wire  \picorv32_core/sel41_b15/B2 ;
  wire  \picorv32_core/sel41_b15/B5 ;
  wire  \picorv32_core/sel41_b16/B2 ;
  wire  \picorv32_core/sel41_b16/B5 ;
  wire  \picorv32_core/sel41_b17/B2 ;
  wire  \picorv32_core/sel41_b17/B5 ;
  wire  \picorv32_core/sel41_b18/B2 ;
  wire  \picorv32_core/sel41_b18/B5 ;
  wire  \picorv32_core/sel41_b19/B2 ;
  wire  \picorv32_core/sel41_b19/B5 ;
  wire  \picorv32_core/sel41_b2/B5 ;
  wire  \picorv32_core/sel41_b20/B2 ;
  wire  \picorv32_core/sel41_b20/B5 ;
  wire  \picorv32_core/sel41_b21/B2 ;
  wire  \picorv32_core/sel41_b21/B5 ;
  wire  \picorv32_core/sel41_b22/B2 ;
  wire  \picorv32_core/sel41_b22/B5 ;
  wire  \picorv32_core/sel41_b23/B2 ;
  wire  \picorv32_core/sel41_b23/B5 ;
  wire  \picorv32_core/sel41_b24/B2 ;
  wire  \picorv32_core/sel41_b24/B5 ;
  wire  \picorv32_core/sel41_b25/B2 ;
  wire  \picorv32_core/sel41_b25/B5 ;
  wire  \picorv32_core/sel41_b26/B2 ;
  wire  \picorv32_core/sel41_b26/B5 ;
  wire  \picorv32_core/sel41_b27/B2 ;
  wire  \picorv32_core/sel41_b27/B5 ;
  wire  \picorv32_core/sel41_b28/B5 ;
  wire  \picorv32_core/sel41_b29/B5 ;
  wire  \picorv32_core/sel41_b3/B5 ;
  wire  \picorv32_core/sel41_b30/B5 ;
  wire  \picorv32_core/sel41_b31/B5 ;
  wire  \picorv32_core/sel41_b4/B2 ;
  wire  \picorv32_core/sel41_b4/B5 ;
  wire  \picorv32_core/sel41_b5/B2 ;
  wire  \picorv32_core/sel41_b5/B5 ;
  wire  \picorv32_core/sel41_b6/B2 ;
  wire  \picorv32_core/sel41_b6/B5 ;
  wire  \picorv32_core/sel41_b7/B2 ;
  wire  \picorv32_core/sel41_b7/B5 ;
  wire  \picorv32_core/sel41_b8/B2 ;
  wire  \picorv32_core/sel41_b8/B5 ;
  wire  \picorv32_core/sel41_b9/B2 ;
  wire  \picorv32_core/sel41_b9/B5 ;
  wire  \picorv32_core/sel42_b0/B4 ;
  wire  \picorv32_core/sel42_b0/B5 ;
  wire  \picorv32_core/sel42_b1/B4 ;
  wire  \picorv32_core/sel42_b1/B5 ;
  wire  \picorv32_core/sel42_b2/B4 ;
  wire  \picorv32_core/sel42_b2/B5 ;
  wire  \picorv32_core/sel42_b3/B4 ;
  wire  \picorv32_core/sel42_b3/B5 ;
  wire  \picorv32_core/sel42_b4/B4 ;
  wire  \picorv32_core/sel42_b4/B5 ;
  wire  \picorv32_core/sel43_b0/B2 ;
  wire  \picorv32_core/sel43_b28/B2 ;
  wire  \picorv32_core/sel43_b29/B2 ;
  wire  \picorv32_core/sel43_b30/B2 ;
  wire  \uart/mux42_b0/B1_1 ;
  wire [3:0] \uart/n35 ;
  wire [3:0] \uart/n4 ;
  wire [3:0] \uart/n49 ;
  wire [31:0] \uart/n5 ;
  wire [3:0] \uart/n50 ;
  wire [4:0] \uart/n57 ;
  wire [3:0] \uart/n77 ;
  wire [31:0] \uart/uart_bsrr ;  // ../src/uart.v(28)
  wire [2:0] \uart/uart_cnt_rx ;  // ../src/uart.v(151)
  wire [31:0] \uart/uart_counter ;  // ../src/uart.v(30)
  wire [7:0] \uart/uart_idr ;  // ../src/uart.v(27)
  wire [7:0] \uart/uart_idr_t ;  // ../src/uart.v(153)
  wire [7:0] \uart/uart_odr ;  // ../src/uart.v(26)
  wire [2:0] \uart/uart_op_clock_by_3_c ;  // ../src/uart.v(35)
  wire [3:0] \uart/uart_smp_rx ;  // ../src/uart.v(152)
  wire [3:0] \uart/uart_status_rxd ;  // ../src/uart.v(148)
  wire [3:0] \uart/uart_status_txd ;  // ../src/uart.v(32)
  wire [31:0] uart_do;  // ../src/top.v(98)
  wire _al_u1001_o;
  wire _al_u1003_o;
  wire _al_u1005_o;
  wire _al_u1007_o;
  wire _al_u1009_o;
  wire _al_u1011_o;
  wire _al_u1013_o;
  wire _al_u1015_o;
  wire _al_u1017_o;
  wire _al_u1019_o;
  wire _al_u1021_o;
  wire _al_u1023_o;
  wire _al_u1025_o;
  wire _al_u1027_o;
  wire _al_u1029_o;
  wire _al_u1031_o;
  wire _al_u1033_o;
  wire _al_u1035_o;
  wire _al_u1037_o;
  wire _al_u1039_o;
  wire _al_u1041_o;
  wire _al_u1043_o;
  wire _al_u1045_o;
  wire _al_u1047_o;
  wire _al_u1049_o;
  wire _al_u1051_o;
  wire _al_u1053_o;
  wire _al_u1055_o;
  wire _al_u1057_o;
  wire _al_u1059_o;
  wire _al_u1061_o;
  wire _al_u1063_o;
  wire _al_u1065_o;
  wire _al_u1066_o;
  wire _al_u1067_o;
  wire _al_u1068_o;
  wire _al_u1070_o;
  wire _al_u1071_o;
  wire _al_u1072_o;
  wire _al_u1074_o;
  wire _al_u1076_o;
  wire _al_u1077_o;
  wire _al_u1079_o;
  wire _al_u1081_o;
  wire _al_u1086_o;
  wire _al_u1088_o;
  wire _al_u1089_o;
  wire _al_u1091_o;
  wire _al_u1092_o;
  wire _al_u1093_o;
  wire _al_u1095_o;
  wire _al_u1096_o;
  wire _al_u1097_o;
  wire _al_u1098_o;
  wire _al_u1100_o;
  wire _al_u1102_o;
  wire _al_u1107_o;
  wire _al_u1108_o;
  wire _al_u1109_o;
  wire _al_u1110_o;
  wire _al_u1111_o;
  wire _al_u1112_o;
  wire _al_u1113_o;
  wire _al_u1117_o;
  wire _al_u1118_o;
  wire _al_u1119_o;
  wire _al_u1120_o;
  wire _al_u1121_o;
  wire _al_u1122_o;
  wire _al_u1123_o;
  wire _al_u1124_o;
  wire _al_u1126_o;
  wire _al_u1127_o;
  wire _al_u1128_o;
  wire _al_u1129_o;
  wire _al_u1130_o;
  wire _al_u1132_o;
  wire _al_u1133_o;
  wire _al_u1134_o;
  wire _al_u1136_o;
  wire _al_u1138_o;
  wire _al_u1140_o;
  wire _al_u1143_o;
  wire _al_u1147_o;
  wire _al_u1151_o;
  wire _al_u1153_o;
  wire _al_u1159_o;
  wire _al_u1160_o;
  wire _al_u1164_o;
  wire _al_u1165_o;
  wire _al_u1168_o;
  wire _al_u1170_o;
  wire _al_u1172_o;
  wire _al_u1173_o;
  wire _al_u1175_o;
  wire _al_u1179_o;
  wire _al_u1183_o;
  wire _al_u1184_o;
  wire _al_u1186_o;
  wire _al_u1187_o;
  wire _al_u1189_o;
  wire _al_u1194_o;
  wire _al_u1195_o;
  wire _al_u1196_o;
  wire _al_u1197_o;
  wire _al_u1198_o;
  wire _al_u1199_o;
  wire _al_u1200_o;
  wire _al_u1201_o;
  wire _al_u1202_o;
  wire _al_u1203_o;
  wire _al_u1204_o;
  wire _al_u1205_o;
  wire _al_u1206_o;
  wire _al_u1207_o;
  wire _al_u1208_o;
  wire _al_u1209_o;
  wire _al_u1210_o;
  wire _al_u1211_o;
  wire _al_u1213_o;
  wire _al_u1214_o;
  wire _al_u1215_o;
  wire _al_u1216_o;
  wire _al_u1218_o;
  wire _al_u1219_o;
  wire _al_u1221_o;
  wire _al_u1224_o;
  wire _al_u1227_o;
  wire _al_u1229_o;
  wire _al_u1230_o;
  wire _al_u1231_o;
  wire _al_u1232_o;
  wire _al_u1235_o;
  wire _al_u1236_o;
  wire _al_u1238_o;
  wire _al_u1239_o;
  wire _al_u1241_o;
  wire _al_u1243_o;
  wire _al_u1245_o;
  wire _al_u1247_o;
  wire _al_u1249_o;
  wire _al_u1251_o;
  wire _al_u1253_o;
  wire _al_u1254_o;
  wire _al_u1257_o;
  wire _al_u1261_o;
  wire _al_u1264_o;
  wire _al_u1266_o;
  wire _al_u1270_o;
  wire _al_u1272_o;
  wire _al_u1273_o;
  wire _al_u1276_o;
  wire _al_u1278_o;
  wire _al_u1279_o;
  wire _al_u1282_o;
  wire _al_u1285_o;
  wire _al_u1288_o;
  wire _al_u1290_o;
  wire _al_u1292_o;
  wire _al_u1293_o;
  wire _al_u1295_o;
  wire _al_u1296_o;
  wire _al_u1298_o;
  wire _al_u1299_o;
  wire _al_u1300_o;
  wire _al_u1301_o;
  wire _al_u1302_o;
  wire _al_u1303_o;
  wire _al_u1304_o;
  wire _al_u1306_o;
  wire _al_u1308_o;
  wire _al_u1310_o;
  wire _al_u1313_o;
  wire _al_u1315_o;
  wire _al_u1319_o;
  wire _al_u1320_o;
  wire _al_u1324_o;
  wire _al_u1325_o;
  wire _al_u1329_o;
  wire _al_u1330_o;
  wire _al_u1334_o;
  wire _al_u1335_o;
  wire _al_u1337_o;
  wire _al_u1338_o;
  wire _al_u1339_o;
  wire _al_u1340_o;
  wire _al_u1343_o;
  wire _al_u1346_o;
  wire _al_u1349_o;
  wire _al_u1352_o;
  wire _al_u1359_o;
  wire _al_u1362_o;
  wire _al_u1367_o;
  wire _al_u1370_o;
  wire _al_u1373_o;
  wire _al_u1376_o;
  wire _al_u1379_o;
  wire _al_u1382_o;
  wire _al_u1385_o;
  wire _al_u1388_o;
  wire _al_u1391_o;
  wire _al_u1394_o;
  wire _al_u1399_o;
  wire _al_u1402_o;
  wire _al_u1405_o;
  wire _al_u1408_o;
  wire _al_u1411_o;
  wire _al_u1414_o;
  wire _al_u1417_o;
  wire _al_u1420_o;
  wire _al_u1423_o;
  wire _al_u1426_o;
  wire _al_u1431_o;
  wire _al_u1432_o;
  wire _al_u1435_o;
  wire _al_u1436_o;
  wire _al_u1439_o;
  wire _al_u1440_o;
  wire _al_u1442_o;
  wire _al_u1443_o;
  wire _al_u1444_o;
  wire _al_u1447_o;
  wire _al_u1448_o;
  wire _al_u1451_o;
  wire _al_u1452_o;
  wire _al_u1456_o;
  wire _al_u1458_o;
  wire _al_u1459_o;
  wire _al_u1464_o;
  wire _al_u1469_o;
  wire _al_u1470_o;
  wire _al_u1481_o;
  wire _al_u1481_o_placeOpt_1;
  wire _al_u1481_o_placeOpt_2;
  wire _al_u1481_o_placeOpt_3;
  wire _al_u1481_o_placeOpt_4;
  wire _al_u1483_o;
  wire _al_u1483_o_placeOpt_1;
  wire _al_u1483_o_placeOpt_2;
  wire _al_u1483_o_placeOpt_3;
  wire _al_u1485_o;
  wire _al_u1485_o_placeOpt_1;
  wire _al_u1485_o_placeOpt_2;
  wire _al_u1485_o_placeOpt_3;
  wire _al_u1493_o;
  wire _al_u1496_o;
  wire _al_u1497_o;
  wire _al_u1498_o;
  wire _al_u1532_o;
  wire _al_u1533_o;
  wire _al_u1535_o;
  wire _al_u1536_o;
  wire _al_u1537_o;
  wire _al_u1538_o;
  wire _al_u1546_o;
  wire _al_u1546_o_placeOpt_1;
  wire _al_u1546_o_placeOpt_2;
  wire _al_u1546_o_placeOpt_3;
  wire _al_u1546_o_placeOpt_4;
  wire _al_u1546_o_placeOpt_5;
  wire _al_u1546_o_placeOpt_6;
  wire _al_u1546_o_placeOpt_7;
  wire _al_u1546_o_placeOpt_8;
  wire _al_u1547_o;
  wire _al_u1548_o;
  wire _al_u1550_o;
  wire _al_u1551_o;
  wire _al_u1552_o;
  wire _al_u1554_o;
  wire _al_u1555_o;
  wire _al_u1557_o;
  wire _al_u1559_o;
  wire _al_u1560_o;
  wire _al_u1563_o;
  wire _al_u1564_o;
  wire _al_u1565_o;
  wire _al_u1566_o;
  wire _al_u1567_o;
  wire _al_u1568_o;
  wire _al_u1569_o;
  wire _al_u1571_o;
  wire _al_u1573_o;
  wire _al_u1575_o;
  wire _al_u1577_o;
  wire _al_u1579_o;
  wire _al_u1580_o;
  wire _al_u1581_o;
  wire _al_u1583_o;
  wire _al_u1585_o;
  wire _al_u1587_o;
  wire _al_u1589_o;
  wire _al_u1591_o;
  wire _al_u1593_o;
  wire _al_u1594_o;
  wire _al_u1596_o;
  wire _al_u1597_o;
  wire _al_u1602_o;
  wire _al_u1603_o;
  wire _al_u1604_o;
  wire _al_u1605_o;
  wire _al_u1606_o;
  wire _al_u1609_o;
  wire _al_u1613_o;
  wire _al_u1614_o;
  wire _al_u1615_o;
  wire _al_u1617_o;
  wire _al_u1618_o;
  wire _al_u1619_o;
  wire _al_u1621_o;
  wire _al_u1622_o;
  wire _al_u1623_o;
  wire _al_u1625_o;
  wire _al_u1626_o;
  wire _al_u1627_o;
  wire _al_u1629_o;
  wire _al_u1630_o;
  wire _al_u1633_o;
  wire _al_u1634_o;
  wire _al_u1635_o;
  wire _al_u1637_o;
  wire _al_u1638_o;
  wire _al_u1640_o;
  wire _al_u1643_o;
  wire _al_u1646_o;
  wire _al_u1648_o;
  wire _al_u1649_o;
  wire _al_u1650_o;
  wire _al_u1651_o;
  wire _al_u1652_o;
  wire _al_u1653_o;
  wire _al_u1654_o;
  wire _al_u1657_o;
  wire _al_u1658_o;
  wire _al_u1660_o;
  wire _al_u1661_o;
  wire _al_u1663_o;
  wire _al_u1664_o;
  wire _al_u1665_o;
  wire _al_u1666_o;
  wire _al_u1667_o;
  wire _al_u1668_o;
  wire _al_u1669_o;
  wire _al_u1672_o;
  wire _al_u1673_o;
  wire _al_u1674_o;
  wire _al_u1675_o;
  wire _al_u1676_o;
  wire _al_u1677_o;
  wire _al_u1679_o;
  wire _al_u1680_o;
  wire _al_u1681_o;
  wire _al_u1682_o;
  wire _al_u1683_o;
  wire _al_u1686_o;
  wire _al_u1687_o;
  wire _al_u1688_o;
  wire _al_u1689_o;
  wire _al_u1690_o;
  wire _al_u1691_o;
  wire _al_u1692_o;
  wire _al_u1695_o;
  wire _al_u1696_o;
  wire _al_u1697_o;
  wire _al_u1698_o;
  wire _al_u1699_o;
  wire _al_u1700_o;
  wire _al_u1701_o;
  wire _al_u1704_o;
  wire _al_u1705_o;
  wire _al_u1706_o;
  wire _al_u1707_o;
  wire _al_u1708_o;
  wire _al_u1709_o;
  wire _al_u1710_o;
  wire _al_u1712_o;
  wire _al_u1713_o;
  wire _al_u1716_o;
  wire _al_u1717_o;
  wire _al_u1718_o;
  wire _al_u1719_o;
  wire _al_u1720_o;
  wire _al_u1723_o;
  wire _al_u1725_o;
  wire _al_u1726_o;
  wire _al_u1727_o;
  wire _al_u1730_o;
  wire _al_u1731_o;
  wire _al_u1734_o;
  wire _al_u1735_o;
  wire _al_u1736_o;
  wire _al_u1737_o;
  wire _al_u1738_o;
  wire _al_u1741_o;
  wire _al_u1743_o;
  wire _al_u1744_o;
  wire _al_u1745_o;
  wire _al_u1748_o;
  wire _al_u1750_o;
  wire _al_u1751_o;
  wire _al_u1752_o;
  wire _al_u1755_o;
  wire _al_u1756_o;
  wire _al_u1757_o;
  wire _al_u1758_o;
  wire _al_u1759_o;
  wire _al_u1762_o;
  wire _al_u1763_o;
  wire _al_u1764_o;
  wire _al_u1765_o;
  wire _al_u1766_o;
  wire _al_u1769_o;
  wire _al_u1770_o;
  wire _al_u1771_o;
  wire _al_u1772_o;
  wire _al_u1773_o;
  wire _al_u1776_o;
  wire _al_u1777_o;
  wire _al_u1778_o;
  wire _al_u1779_o;
  wire _al_u1780_o;
  wire _al_u1783_o;
  wire _al_u1784_o;
  wire _al_u1785_o;
  wire _al_u1786_o;
  wire _al_u1787_o;
  wire _al_u1790_o;
  wire _al_u1791_o;
  wire _al_u1792_o;
  wire _al_u1793_o;
  wire _al_u1794_o;
  wire _al_u1797_o;
  wire _al_u1798_o;
  wire _al_u1799_o;
  wire _al_u1800_o;
  wire _al_u1801_o;
  wire _al_u1804_o;
  wire _al_u1805_o;
  wire _al_u1806_o;
  wire _al_u1807_o;
  wire _al_u1808_o;
  wire _al_u1811_o;
  wire _al_u1812_o;
  wire _al_u1814_o;
  wire _al_u1815_o;
  wire _al_u1816_o;
  wire _al_u1817_o;
  wire _al_u1818_o;
  wire _al_u1821_o;
  wire _al_u1822_o;
  wire _al_u1823_o;
  wire _al_u1824_o;
  wire _al_u1825_o;
  wire _al_u1828_o;
  wire _al_u1829_o;
  wire _al_u1830_o;
  wire _al_u1831_o;
  wire _al_u1832_o;
  wire _al_u1835_o;
  wire _al_u1836_o;
  wire _al_u1837_o;
  wire _al_u1838_o;
  wire _al_u1839_o;
  wire _al_u1842_o;
  wire _al_u1843_o;
  wire _al_u1844_o;
  wire _al_u1845_o;
  wire _al_u1846_o;
  wire _al_u1848_o;
  wire _al_u1849_o;
  wire _al_u1850_o;
  wire _al_u1851_o;
  wire _al_u1852_o;
  wire _al_u1853_o;
  wire _al_u1855_o;
  wire _al_u1856_o;
  wire _al_u1857_o;
  wire _al_u1858_o;
  wire _al_u1859_o;
  wire _al_u1860_o;
  wire _al_u1862_o;
  wire _al_u1863_o;
  wire _al_u1864_o;
  wire _al_u1865_o;
  wire _al_u1866_o;
  wire _al_u1867_o;
  wire _al_u1869_o;
  wire _al_u1870_o;
  wire _al_u1871_o;
  wire _al_u1872_o;
  wire _al_u1873_o;
  wire _al_u1874_o;
  wire _al_u1876_o;
  wire _al_u1877_o;
  wire _al_u1878_o;
  wire _al_u1879_o;
  wire _al_u1880_o;
  wire _al_u1881_o;
  wire _al_u1883_o;
  wire _al_u1884_o;
  wire _al_u1885_o;
  wire _al_u1886_o;
  wire _al_u1887_o;
  wire _al_u1888_o;
  wire _al_u1890_o;
  wire _al_u1891_o;
  wire _al_u1892_o;
  wire _al_u1893_o;
  wire _al_u1894_o;
  wire _al_u1895_o;
  wire _al_u1898_o;
  wire _al_u1899_o;
  wire _al_u1900_o;
  wire _al_u1902_o;
  wire _al_u1903_o;
  wire _al_u1904_o;
  wire _al_u1906_o;
  wire _al_u1908_o;
  wire _al_u1909_o;
  wire _al_u1910_o;
  wire _al_u1911_o;
  wire _al_u1912_o;
  wire _al_u1914_o;
  wire _al_u1915_o;
  wire _al_u1916_o;
  wire _al_u1917_o;
  wire _al_u1918_o;
  wire _al_u1920_o;
  wire _al_u1921_o;
  wire _al_u1922_o;
  wire _al_u1923_o;
  wire _al_u1924_o;
  wire _al_u1925_o;
  wire _al_u1926_o;
  wire _al_u1927_o;
  wire _al_u1929_o;
  wire _al_u1930_o;
  wire _al_u1932_o;
  wire _al_u1934_o;
  wire _al_u1935_o;
  wire _al_u1936_o;
  wire _al_u1937_o;
  wire _al_u1938_o;
  wire _al_u1940_o;
  wire _al_u1941_o;
  wire _al_u1943_o;
  wire _al_u1945_o;
  wire _al_u1946_o;
  wire _al_u1947_o;
  wire _al_u1948_o;
  wire _al_u1949_o;
  wire _al_u1951_o;
  wire _al_u1952_o;
  wire _al_u1954_o;
  wire _al_u1956_o;
  wire _al_u1957_o;
  wire _al_u1958_o;
  wire _al_u1959_o;
  wire _al_u1960_o;
  wire _al_u1962_o;
  wire _al_u1963_o;
  wire _al_u1965_o;
  wire _al_u1967_o;
  wire _al_u1968_o;
  wire _al_u1969_o;
  wire _al_u1970_o;
  wire _al_u1971_o;
  wire _al_u1973_o;
  wire _al_u1974_o;
  wire _al_u1976_o;
  wire _al_u1978_o;
  wire _al_u1979_o;
  wire _al_u1980_o;
  wire _al_u1981_o;
  wire _al_u1982_o;
  wire _al_u1984_o;
  wire _al_u1985_o;
  wire _al_u1987_o;
  wire _al_u1989_o;
  wire _al_u1990_o;
  wire _al_u1991_o;
  wire _al_u1992_o;
  wire _al_u1993_o;
  wire _al_u1995_o;
  wire _al_u1996_o;
  wire _al_u1997_o;
  wire _al_u1999_o;
  wire _al_u2000_o;
  wire _al_u2001_o;
  wire _al_u2002_o;
  wire _al_u2003_o;
  wire _al_u2005_o;
  wire _al_u2007_o;
  wire _al_u2009_o;
  wire _al_u2010_o;
  wire _al_u2011_o;
  wire _al_u2012_o;
  wire _al_u2013_o;
  wire _al_u2014_o;
  wire _al_u2015_o;
  wire _al_u2016_o;
  wire _al_u2018_o;
  wire _al_u2020_o;
  wire _al_u2021_o;
  wire _al_u2022_o;
  wire _al_u2023_o;
  wire _al_u2024_o;
  wire _al_u2026_o;
  wire _al_u2027_o;
  wire _al_u2028_o;
  wire _al_u2030_o;
  wire _al_u2031_o;
  wire _al_u2032_o;
  wire _al_u2033_o;
  wire _al_u2034_o;
  wire _al_u2035_o;
  wire _al_u2036_o;
  wire _al_u2038_o;
  wire _al_u2040_o;
  wire _al_u2041_o;
  wire _al_u2042_o;
  wire _al_u2043_o;
  wire _al_u2044_o;
  wire _al_u2045_o;
  wire _al_u2046_o;
  wire _al_u2048_o;
  wire _al_u2050_o;
  wire _al_u2051_o;
  wire _al_u2052_o;
  wire _al_u2053_o;
  wire _al_u2054_o;
  wire _al_u2056_o;
  wire _al_u2057_o;
  wire _al_u2059_o;
  wire _al_u2061_o;
  wire _al_u2062_o;
  wire _al_u2063_o;
  wire _al_u2064_o;
  wire _al_u2065_o;
  wire _al_u2067_o;
  wire _al_u2068_o;
  wire _al_u2070_o;
  wire _al_u2072_o;
  wire _al_u2073_o;
  wire _al_u2074_o;
  wire _al_u2075_o;
  wire _al_u2076_o;
  wire _al_u2078_o;
  wire _al_u2079_o;
  wire _al_u2081_o;
  wire _al_u2083_o;
  wire _al_u2084_o;
  wire _al_u2085_o;
  wire _al_u2086_o;
  wire _al_u2087_o;
  wire _al_u2089_o;
  wire _al_u2090_o;
  wire _al_u2092_o;
  wire _al_u2094_o;
  wire _al_u2095_o;
  wire _al_u2096_o;
  wire _al_u2097_o;
  wire _al_u2098_o;
  wire _al_u2100_o;
  wire _al_u2101_o;
  wire _al_u2103_o;
  wire _al_u2105_o;
  wire _al_u2106_o;
  wire _al_u2107_o;
  wire _al_u2108_o;
  wire _al_u2109_o;
  wire _al_u2111_o;
  wire _al_u2112_o;
  wire _al_u2114_o;
  wire _al_u2116_o;
  wire _al_u2117_o;
  wire _al_u2118_o;
  wire _al_u2119_o;
  wire _al_u2120_o;
  wire _al_u2122_o;
  wire _al_u2123_o;
  wire _al_u2125_o;
  wire _al_u2127_o;
  wire _al_u2128_o;
  wire _al_u2129_o;
  wire _al_u2130_o;
  wire _al_u2131_o;
  wire _al_u2133_o;
  wire _al_u2134_o;
  wire _al_u2136_o;
  wire _al_u2138_o;
  wire _al_u2139_o;
  wire _al_u2140_o;
  wire _al_u2141_o;
  wire _al_u2142_o;
  wire _al_u2144_o;
  wire _al_u2145_o;
  wire _al_u2146_o;
  wire _al_u2148_o;
  wire _al_u2149_o;
  wire _al_u2150_o;
  wire _al_u2151_o;
  wire _al_u2152_o;
  wire _al_u2154_o;
  wire _al_u2155_o;
  wire _al_u2157_o;
  wire _al_u2159_o;
  wire _al_u2160_o;
  wire _al_u2161_o;
  wire _al_u2162_o;
  wire _al_u2163_o;
  wire _al_u2165_o;
  wire _al_u2166_o;
  wire _al_u2168_o;
  wire _al_u2170_o;
  wire _al_u2171_o;
  wire _al_u2172_o;
  wire _al_u2173_o;
  wire _al_u2174_o;
  wire _al_u2176_o;
  wire _al_u2177_o;
  wire _al_u2179_o;
  wire _al_u2181_o;
  wire _al_u2182_o;
  wire _al_u2183_o;
  wire _al_u2184_o;
  wire _al_u2185_o;
  wire _al_u2187_o;
  wire _al_u2188_o;
  wire _al_u2190_o;
  wire _al_u2192_o;
  wire _al_u2193_o;
  wire _al_u2194_o;
  wire _al_u2195_o;
  wire _al_u2196_o;
  wire _al_u2198_o;
  wire _al_u2199_o;
  wire _al_u2201_o;
  wire _al_u2203_o;
  wire _al_u2204_o;
  wire _al_u2205_o;
  wire _al_u2206_o;
  wire _al_u2207_o;
  wire _al_u2209_o;
  wire _al_u2210_o;
  wire _al_u2212_o;
  wire _al_u2214_o;
  wire _al_u2215_o;
  wire _al_u2216_o;
  wire _al_u2217_o;
  wire _al_u2218_o;
  wire _al_u2220_o;
  wire _al_u2221_o;
  wire _al_u2223_o;
  wire _al_u2225_o;
  wire _al_u2226_o;
  wire _al_u2227_o;
  wire _al_u2228_o;
  wire _al_u2229_o;
  wire _al_u2231_o;
  wire _al_u2232_o;
  wire _al_u2234_o;
  wire _al_u2236_o;
  wire _al_u2237_o;
  wire _al_u2238_o;
  wire _al_u2239_o;
  wire _al_u2240_o;
  wire _al_u2242_o;
  wire _al_u2243_o;
  wire _al_u2245_o;
  wire _al_u2247_o;
  wire _al_u2248_o;
  wire _al_u2249_o;
  wire _al_u2250_o;
  wire _al_u2251_o;
  wire _al_u2253_o;
  wire _al_u2254_o;
  wire _al_u2256_o;
  wire _al_u2258_o;
  wire _al_u2259_o;
  wire _al_u2260_o;
  wire _al_u2261_o;
  wire _al_u2262_o;
  wire _al_u2263_o;
  wire _al_u2265_o;
  wire _al_u2267_o;
  wire _al_u2268_o;
  wire _al_u2269_o;
  wire _al_u2270_o;
  wire _al_u2271_o;
  wire _al_u2272_o;
  wire _al_u2273_o;
  wire _al_u2274_o;
  wire _al_u2275_o;
  wire _al_u2276_o;
  wire _al_u2277_o;
  wire _al_u2278_o;
  wire _al_u2279_o;
  wire _al_u2281_o;
  wire _al_u2282_o;
  wire _al_u2283_o;
  wire _al_u2284_o;
  wire _al_u2285_o;
  wire _al_u2287_o;
  wire _al_u2288_o;
  wire _al_u2289_o;
  wire _al_u2290_o;
  wire _al_u2291_o;
  wire _al_u2292_o;
  wire _al_u2293_o;
  wire _al_u2294_o;
  wire _al_u2295_o;
  wire _al_u2296_o;
  wire _al_u2297_o;
  wire _al_u2301_o;
  wire _al_u2302_o;
  wire _al_u2305_o;
  wire _al_u2306_o;
  wire _al_u2307_o;
  wire _al_u2309_o;
  wire _al_u2310_o;
  wire _al_u2315_o;
  wire _al_u2316_o;
  wire _al_u2317_o;
  wire _al_u2318_o;
  wire _al_u2319_o;
  wire _al_u2320_o;
  wire _al_u2321_o;
  wire _al_u2322_o;
  wire _al_u2323_o;
  wire _al_u2324_o;
  wire _al_u2325_o;
  wire _al_u2327_o;
  wire _al_u2328_o;
  wire _al_u2329_o;
  wire _al_u2330_o;
  wire _al_u2331_o;
  wire _al_u2332_o;
  wire _al_u2333_o;
  wire _al_u2334_o;
  wire _al_u2335_o;
  wire _al_u2337_o;
  wire _al_u2338_o;
  wire _al_u2339_o;
  wire _al_u2340_o;
  wire _al_u2341_o;
  wire _al_u2342_o;
  wire _al_u2344_o;
  wire _al_u2345_o;
  wire _al_u2346_o;
  wire _al_u2347_o;
  wire _al_u2348_o;
  wire _al_u2349_o;
  wire _al_u2350_o;
  wire _al_u2351_o;
  wire _al_u2353_o;
  wire _al_u2354_o;
  wire _al_u2355_o;
  wire _al_u2356_o;
  wire _al_u2357_o;
  wire _al_u2358_o;
  wire _al_u2359_o;
  wire _al_u2360_o;
  wire _al_u2363_o;
  wire _al_u2364_o;
  wire _al_u2365_o;
  wire _al_u2366_o;
  wire _al_u2367_o;
  wire _al_u2368_o;
  wire _al_u2370_o;
  wire _al_u2371_o;
  wire _al_u2372_o;
  wire _al_u2373_o;
  wire _al_u2374_o;
  wire _al_u2375_o;
  wire _al_u2376_o;
  wire _al_u2377_o;
  wire _al_u2378_o;
  wire _al_u2379_o;
  wire _al_u2380_o;
  wire _al_u2382_o;
  wire _al_u2383_o;
  wire _al_u2384_o;
  wire _al_u2385_o;
  wire _al_u2386_o;
  wire _al_u2387_o;
  wire _al_u2388_o;
  wire _al_u2389_o;
  wire _al_u2390_o;
  wire _al_u2391_o;
  wire _al_u2392_o;
  wire _al_u2393_o;
  wire _al_u2395_o;
  wire _al_u2396_o;
  wire _al_u2397_o;
  wire _al_u2398_o;
  wire _al_u2399_o;
  wire _al_u2400_o;
  wire _al_u2401_o;
  wire _al_u2402_o;
  wire _al_u2403_o;
  wire _al_u2404_o;
  wire _al_u2405_o;
  wire _al_u2406_o;
  wire _al_u2408_o;
  wire _al_u2410_o;
  wire _al_u2411_o;
  wire _al_u2412_o;
  wire _al_u2413_o;
  wire _al_u2414_o;
  wire _al_u2415_o;
  wire _al_u2416_o;
  wire _al_u2417_o;
  wire _al_u2418_o;
  wire _al_u2420_o;
  wire _al_u2421_o;
  wire _al_u2422_o;
  wire _al_u2424_o;
  wire _al_u2425_o;
  wire _al_u2426_o;
  wire _al_u2427_o;
  wire _al_u2429_o;
  wire _al_u2430_o;
  wire _al_u2431_o;
  wire _al_u2433_o;
  wire _al_u2434_o;
  wire _al_u2435_o;
  wire _al_u2436_o;
  wire _al_u2437_o;
  wire _al_u2440_o;
  wire _al_u2441_o;
  wire _al_u2443_o;
  wire _al_u2444_o;
  wire _al_u2446_o;
  wire _al_u2447_o;
  wire _al_u2449_o;
  wire _al_u2450_o;
  wire _al_u2451_o;
  wire _al_u2453_o;
  wire _al_u2454_o;
  wire _al_u2455_o;
  wire _al_u2457_o;
  wire _al_u2458_o;
  wire _al_u2459_o;
  wire _al_u2460_o;
  wire _al_u2461_o;
  wire _al_u2462_o;
  wire _al_u2464_o;
  wire _al_u2465_o;
  wire _al_u2466_o;
  wire _al_u2467_o;
  wire _al_u2468_o;
  wire _al_u2469_o;
  wire _al_u2470_o;
  wire _al_u2471_o;
  wire _al_u2473_o;
  wire _al_u2474_o;
  wire _al_u2475_o;
  wire _al_u2476_o;
  wire _al_u2477_o;
  wire _al_u2478_o;
  wire _al_u2479_o;
  wire _al_u665_o;
  wire _al_u700_o;
  wire _al_u700_o_placeOpt_1;
  wire _al_u700_o_placeOpt_2;
  wire _al_u700_o_placeOpt_3;
  wire _al_u799_o;
  wire _al_u803_o;
  wire _al_u810_o;
  wire _al_u811_o;
  wire _al_u812_o;
  wire _al_u813_o;
  wire _al_u815_o;
  wire _al_u816_o;
  wire _al_u817_o;
  wire _al_u826_o;
  wire _al_u827_o;
  wire _al_u828_o;
  wire _al_u829_o;
  wire _al_u831_o;
  wire _al_u833_o;
  wire _al_u835_o;
  wire _al_u837_o;
  wire _al_u839_o;
  wire _al_u841_o;
  wire _al_u843_o;
  wire _al_u845_o;
  wire _al_u847_o;
  wire _al_u849_o;
  wire _al_u851_o;
  wire _al_u853_o;
  wire _al_u855_o;
  wire _al_u857_o;
  wire _al_u859_o;
  wire _al_u861_o;
  wire _al_u863_o;
  wire _al_u865_o;
  wire _al_u867_o;
  wire _al_u869_o;
  wire _al_u871_o;
  wire _al_u873_o;
  wire _al_u875_o;
  wire _al_u877_o;
  wire _al_u879_o;
  wire _al_u881_o;
  wire _al_u883_o;
  wire _al_u885_o;
  wire _al_u887_o;
  wire _al_u889_o;
  wire _al_u892_o;
  wire _al_u893_o;
  wire _al_u894_o;
  wire _al_u896_o;
  wire _al_u902_o;
  wire _al_u904_o;
  wire _al_u906_o;
  wire _al_u908_o;
  wire _al_u909_o;
  wire _al_u930_o;
  wire _al_u933_o;
  wire _al_u973_o;
  wire _al_u976_o;
  wire _al_u979_o;
  wire _al_u980_o;
  wire _al_u982_o;
  wire _al_u999_o;
  wire clk_pad;  // ../src/top.v(4)
  wire \eq0/or_xor_i0$0$_i1$0$_o_o ;
  wire \eq1/or_xor_i0$13$_i1$13$_o_lutinv ;
  wire \eq1/or_xor_i0$17$_i1$17$_o_lutinv ;
  wire \eq2/or_xor_i0$1$_i1$1$_o_o_lutinv ;
  wire \eq2/or_xor_i0$5$_i1$5$_o_o_lutinv ;
  wire n11;
  wire n13;
  wire n16;
  wire n7;
  wire n9;
  wire \picorv32_core/add0/c1 ;
  wire \picorv32_core/add0/c11 ;
  wire \picorv32_core/add0/c13 ;
  wire \picorv32_core/add0/c15 ;
  wire \picorv32_core/add0/c17 ;
  wire \picorv32_core/add0/c19 ;
  wire \picorv32_core/add0/c21 ;
  wire \picorv32_core/add0/c23 ;
  wire \picorv32_core/add0/c25 ;
  wire \picorv32_core/add0/c27 ;
  wire \picorv32_core/add0/c29 ;
  wire \picorv32_core/add0/c3 ;
  wire \picorv32_core/add0/c5 ;
  wire \picorv32_core/add0/c7 ;
  wire \picorv32_core/add0/c9 ;
  wire \picorv32_core/add1/c11 ;
  wire \picorv32_core/add1/c15 ;
  wire \picorv32_core/add1/c19 ;
  wire \picorv32_core/add1/c23 ;
  wire \picorv32_core/add1/c27 ;
  wire \picorv32_core/add1/c3 ;
  wire \picorv32_core/add1/c31 ;
  wire \picorv32_core/add1/c7 ;
  wire \picorv32_core/add2/c11 ;
  wire \picorv32_core/add2/c15 ;
  wire \picorv32_core/add2/c19 ;
  wire \picorv32_core/add2/c23 ;
  wire \picorv32_core/add2/c27 ;
  wire \picorv32_core/add2/c3 ;
  wire \picorv32_core/add2/c31 ;
  wire \picorv32_core/add2/c7 ;
  wire \picorv32_core/add3/c11 ;
  wire \picorv32_core/add3/c15 ;
  wire \picorv32_core/add3/c19 ;
  wire \picorv32_core/add3/c23 ;
  wire \picorv32_core/add3/c27 ;
  wire \picorv32_core/add3/c3 ;
  wire \picorv32_core/add3/c31 ;
  wire \picorv32_core/add3/c35 ;
  wire \picorv32_core/add3/c39 ;
  wire \picorv32_core/add3/c43 ;
  wire \picorv32_core/add3/c47 ;
  wire \picorv32_core/add3/c51 ;
  wire \picorv32_core/add3/c55 ;
  wire \picorv32_core/add3/c59 ;
  wire \picorv32_core/add3/c63 ;
  wire \picorv32_core/add3/c7 ;
  wire \picorv32_core/add4/c11 ;
  wire \picorv32_core/add4/c15 ;
  wire \picorv32_core/add4/c19 ;
  wire \picorv32_core/add4/c23 ;
  wire \picorv32_core/add4/c27 ;
  wire \picorv32_core/add4/c3 ;
  wire \picorv32_core/add4/c31 ;
  wire \picorv32_core/add4/c7 ;
  wire \picorv32_core/add5/c11 ;
  wire \picorv32_core/add5/c15 ;
  wire \picorv32_core/add5/c19 ;
  wire \picorv32_core/add5/c23 ;
  wire \picorv32_core/add5/c27 ;
  wire \picorv32_core/add5/c3 ;
  wire \picorv32_core/add5/c31 ;
  wire \picorv32_core/add5/c35 ;
  wire \picorv32_core/add5/c39 ;
  wire \picorv32_core/add5/c43 ;
  wire \picorv32_core/add5/c47 ;
  wire \picorv32_core/add5/c51 ;
  wire \picorv32_core/add5/c55 ;
  wire \picorv32_core/add5/c59 ;
  wire \picorv32_core/add5/c63 ;
  wire \picorv32_core/add5/c7 ;
  wire \picorv32_core/add6/c11 ;
  wire \picorv32_core/add6/c15 ;
  wire \picorv32_core/add6/c19 ;
  wire \picorv32_core/add6/c23 ;
  wire \picorv32_core/add6/c27 ;
  wire \picorv32_core/add6/c3 ;
  wire \picorv32_core/add6/c31 ;
  wire \picorv32_core/add6/c7 ;
  wire \picorv32_core/add7/c11 ;
  wire \picorv32_core/add7/c15 ;
  wire \picorv32_core/add7/c19 ;
  wire \picorv32_core/add7/c23 ;
  wire \picorv32_core/add7/c27 ;
  wire \picorv32_core/add7/c3 ;
  wire \picorv32_core/add7/c31 ;
  wire \picorv32_core/add7/c7 ;
  wire \picorv32_core/add8/c1 ;
  wire \picorv32_core/add8/c11 ;
  wire \picorv32_core/add8/c13 ;
  wire \picorv32_core/add8/c15 ;
  wire \picorv32_core/add8/c17 ;
  wire \picorv32_core/add8/c19 ;
  wire \picorv32_core/add8/c21 ;
  wire \picorv32_core/add8/c23 ;
  wire \picorv32_core/add8/c25 ;
  wire \picorv32_core/add8/c27 ;
  wire \picorv32_core/add8/c29 ;
  wire \picorv32_core/add8/c3 ;
  wire \picorv32_core/add8/c31 ;
  wire \picorv32_core/add8/c5 ;
  wire \picorv32_core/add8/c7 ;
  wire \picorv32_core/add8/c9 ;
  wire \picorv32_core/alu_eq_lutinv ;  // ../src/picorv32.v(1180)
  wire \picorv32_core/alu_lts ;  // ../src/picorv32.v(1180)
  wire \picorv32_core/alu_ltu ;  // ../src/picorv32.v(1180)
  wire \picorv32_core/clear_prefetched_high_word_q ;  // ../src/picorv32.v(1240)
  wire \picorv32_core/compressed_instr ;  // ../src/picorv32.v(625)
  wire \picorv32_core/cpuregs_p1/dram_do_i0_000 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_001 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_002 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_003 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_004 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_005 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_006 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_007 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_008 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_009 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_010 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_011 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_012 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_013 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_014 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_015 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_016 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_017 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_018 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_019 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_020 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_021 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_022 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_023 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_024 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_025 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_026 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_027 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_028 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_029 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_030 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i0_031 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_000 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_001 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_002 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_003 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_004 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_005 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_006 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_007 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_008 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_009 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_010 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_011 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_012 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_013 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_014 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_015 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_016 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_017 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_018 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_019 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_020 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_021 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_022 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_023 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_024 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_025 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_026 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_027 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_028 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_029 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_030 ;
  wire \picorv32_core/cpuregs_p1/dram_do_i1_031 ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c0_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c0_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c0_we ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c1_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c1_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c1_we ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c2_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c2_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c2_we ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c3_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c3_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c3_we ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c4_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c4_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c4_we ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c5_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c5_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c5_we ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c6_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c6_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c6_we ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c7_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c7_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r0_c7_we ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c0_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c0_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c0_we ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c1_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c1_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c1_we ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c2_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c2_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c2_we ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c3_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c3_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c3_we ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c4_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c4_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c4_we ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c5_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c5_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c5_we ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c6_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c6_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c6_we ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c7_mode ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c7_wclk ;
  wire \picorv32_core/cpuregs_p1/dram_r1_c7_we ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_000 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_001 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_002 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_003 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_004 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_005 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_006 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_007 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_008 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_009 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_010 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_011 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_012 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_013 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_014 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_015 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_016 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_017 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_018 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_019 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_020 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_021 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_022 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_023 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_024 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_025 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_026 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_027 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_028 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_029 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_030 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i0_031 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_000 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_001 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_002 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_003 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_004 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_005 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_006 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_007 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_008 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_009 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_010 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_011 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_012 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_013 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_014 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_015 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_016 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_017 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_018 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_019 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_020 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_021 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_022 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_023 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_024 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_025 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_026 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_027 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_028 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_029 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_030 ;
  wire \picorv32_core/cpuregs_p2/dram_do_i1_031 ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c0_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c0_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c0_we ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c1_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c1_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c1_we ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c2_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c2_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c2_we ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c3_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c3_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c3_we ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c4_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c4_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c4_we ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c5_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c5_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c5_we ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c6_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c6_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c6_we ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c7_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c7_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r0_c7_we ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c0_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c0_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c0_we ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c1_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c1_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c1_we ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c2_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c2_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c2_we ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c3_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c3_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c3_we ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c4_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c4_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c4_we ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c5_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c5_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c5_we ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c6_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c6_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c6_we ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c7_mode ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c7_wclk ;
  wire \picorv32_core/cpuregs_p2/dram_r1_c7_we ;
  wire \picorv32_core/decoder_pseudo_trigger ;  // ../src/picorv32.v(623)
  wire \picorv32_core/decoder_trigger ;  // ../src/picorv32.v(621)
  wire \picorv32_core/instr_add ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_addi ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_and ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_andi ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_auipc ;  // ../src/picorv32.v(610)
  wire \picorv32_core/instr_beq ;  // ../src/picorv32.v(611)
  wire \picorv32_core/instr_bge ;  // ../src/picorv32.v(611)
  wire \picorv32_core/instr_bgeu ;  // ../src/picorv32.v(611)
  wire \picorv32_core/instr_blt ;  // ../src/picorv32.v(611)
  wire \picorv32_core/instr_bltu ;  // ../src/picorv32.v(611)
  wire \picorv32_core/instr_bne ;  // ../src/picorv32.v(611)
  wire \picorv32_core/instr_jal ;  // ../src/picorv32.v(610)
  wire \picorv32_core/instr_jalr ;  // ../src/picorv32.v(610)
  wire \picorv32_core/instr_lb ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_lbu ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_lh ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_lhu ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_lui ;  // ../src/picorv32.v(610)
  wire \picorv32_core/instr_lw ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_or ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_ori ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_rdcycle ;  // ../src/picorv32.v(615)
  wire \picorv32_core/instr_rdcycleh ;  // ../src/picorv32.v(615)
  wire \picorv32_core/instr_rdinstr ;  // ../src/picorv32.v(615)
  wire \picorv32_core/instr_rdinstrh ;  // ../src/picorv32.v(615)
  wire \picorv32_core/instr_sb ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_sh ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_sll ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_slli ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_slt ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_slti ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_sltiu ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_sltu ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_sra ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_srai ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_srl ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_srli ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_sub ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_sw ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_xor ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_xori ;  // ../src/picorv32.v(613)
  wire \picorv32_core/is_alu_reg_imm ;  // ../src/picorv32.v(638)
  wire \picorv32_core/is_alu_reg_reg ;  // ../src/picorv32.v(639)
  wire \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ;  // ../src/picorv32.v(636)
  wire \picorv32_core/is_compare ;  // ../src/picorv32.v(640)
  wire \picorv32_core/is_jalr_addi_slti_sltiu_xori_ori_andi ;  // ../src/picorv32.v(630)
  wire \picorv32_core/is_lb_lh_lw_lbu_lhu ;  // ../src/picorv32.v(628)
  wire \picorv32_core/is_lbu_lhu_lw ;  // ../src/picorv32.v(637)
  wire \picorv32_core/is_lui_auipc_jal ;  // ../src/picorv32.v(627)
  wire \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub ;  // ../src/picorv32.v(633)
  wire \picorv32_core/is_sb_sh_sw ;  // ../src/picorv32.v(631)
  wire \picorv32_core/is_sll_srl_sra ;  // ../src/picorv32.v(632)
  wire \picorv32_core/is_slli_srli_srai ;  // ../src/picorv32.v(629)
  wire \picorv32_core/is_slti_blt_slt ;  // ../src/picorv32.v(634)
  wire \picorv32_core/is_sltiu_bltu_sltu ;  // ../src/picorv32.v(635)
  wire \picorv32_core/latched_branch ;  // ../src/picorv32.v(1157)
  wire \picorv32_core/latched_compr ;  // ../src/picorv32.v(1158)
  wire \picorv32_core/latched_is_lb ;  // ../src/picorv32.v(1162)
  wire \picorv32_core/latched_is_lh ;  // ../src/picorv32.v(1161)
  wire \picorv32_core/latched_is_lu ;  // ../src/picorv32.v(1160)
  wire \picorv32_core/latched_stalu ;  // ../src/picorv32.v(1156)
  wire \picorv32_core/latched_store ;  // ../src/picorv32.v(1155)
  wire \picorv32_core/lt0_c1 ;
  wire \picorv32_core/lt0_c11 ;
  wire \picorv32_core/lt0_c13 ;
  wire \picorv32_core/lt0_c15 ;
  wire \picorv32_core/lt0_c17 ;
  wire \picorv32_core/lt0_c19 ;
  wire \picorv32_core/lt0_c21 ;
  wire \picorv32_core/lt0_c23 ;
  wire \picorv32_core/lt0_c25 ;
  wire \picorv32_core/lt0_c27 ;
  wire \picorv32_core/lt0_c29 ;
  wire \picorv32_core/lt0_c3 ;
  wire \picorv32_core/lt0_c31 ;
  wire \picorv32_core/lt0_c5 ;
  wire \picorv32_core/lt0_c7 ;
  wire \picorv32_core/lt0_c9 ;
  wire \picorv32_core/lt1_c1 ;
  wire \picorv32_core/lt1_c11 ;
  wire \picorv32_core/lt1_c13 ;
  wire \picorv32_core/lt1_c15 ;
  wire \picorv32_core/lt1_c17 ;
  wire \picorv32_core/lt1_c19 ;
  wire \picorv32_core/lt1_c21 ;
  wire \picorv32_core/lt1_c23 ;
  wire \picorv32_core/lt1_c25 ;
  wire \picorv32_core/lt1_c27 ;
  wire \picorv32_core/lt1_c29 ;
  wire \picorv32_core/lt1_c3 ;
  wire \picorv32_core/lt1_c31 ;
  wire \picorv32_core/lt1_c5 ;
  wire \picorv32_core/lt1_c7 ;
  wire \picorv32_core/lt1_c9 ;
  wire \picorv32_core/lt2_c1 ;
  wire \picorv32_core/lt2_c3 ;
  wire \picorv32_core/lt2_c5 ;
  wire \picorv32_core/mem_do_prefetch ;  // ../src/picorv32.v(320)
  wire \picorv32_core/mem_do_prefetch_placeOpt_1 ;
  wire \picorv32_core/mem_do_prefetch_placeOpt_2 ;
  wire \picorv32_core/mem_do_prefetch_placeOpt_3 ;
  wire \picorv32_core/mem_do_prefetch_placeOpt_4 ;
  wire \picorv32_core/mem_do_prefetch_placeOpt_5 ;
  wire \picorv32_core/mem_do_prefetch_placeOpt_6 ;
  wire \picorv32_core/mem_do_prefetch_placeOpt_7 ;
  wire \picorv32_core/mem_do_prefetch_placeOpt_8 ;
  wire \picorv32_core/mem_do_rdata ;  // ../src/picorv32.v(322)
  wire \picorv32_core/mem_do_rinst ;  // ../src/picorv32.v(321)
  wire \picorv32_core/mem_do_wdata ;  // ../src/picorv32.v(323)
  wire \picorv32_core/mem_la_firstword_xfer ;  // ../src/picorv32.v(327)
  wire \picorv32_core/mem_la_read ;  // ../src/picorv32.v(87)
  wire \picorv32_core/mem_la_secondword ;  // ../src/picorv32.v(325)
  wire \picorv32_core/mem_rdata_latched$0$_placeOpt_1 ;
  wire \picorv32_core/mem_rdata_latched$0$_placeOpt_2 ;
  wire \picorv32_core/mem_rdata_latched$0$_placeOpt_3 ;
  wire \picorv32_core/mem_rdata_latched$0$_placeOpt_4 ;
  wire \picorv32_core/mem_rdata_latched$0$_placeOpt_5 ;
  wire \picorv32_core/mem_rdata_latched$1$_placeOpt_1 ;
  wire \picorv32_core/mem_rdata_latched$1$_placeOpt_2 ;
  wire \picorv32_core/mem_rdata_latched$1$_placeOpt_3 ;
  wire \picorv32_core/mem_rdata_latched$1$_placeOpt_4 ;
  wire \picorv32_core/mem_valid ;  // ../src/picorv32.v(77)
  wire \picorv32_core/mem_xfer ;  // ../src/picorv32.v(337)
  wire \picorv32_core/mem_xfer_placeOpt_1 ;
  wire \picorv32_core/mem_xfer_placeOpt_2 ;
  wire \picorv32_core/mem_xfer_placeOpt_3 ;
  wire \picorv32_core/mem_xfer_placeOpt_4 ;
  wire \picorv32_core/mem_xfer_placeOpt_5 ;
  wire \picorv32_core/mux132_b0_sel_is_3_o ;
  wire \picorv32_core/mux164_b0_sel_is_0_o ;
  wire \picorv32_core/mux3_b16_sel_is_0_o ;
  wire \picorv32_core/mux4_b0_sel_is_0_o ;
  wire \picorv32_core/mux51_b0_sel_is_3_o ;
  wire \picorv32_core/mux59_sel_is_5_o ;
  wire \picorv32_core/mux61_sel_is_5_o ;
  wire \picorv32_core/mux68_b0_sel_is_2_o ;
  wire \picorv32_core/mux81_sel_is_1_o ;
  wire \picorv32_core/n111 ;
  wire \picorv32_core/n131 ;
  wire \picorv32_core/n15_lutinv ;
  wire \picorv32_core/n16 ;
  wire \picorv32_core/n165 ;
  wire \picorv32_core/n168 ;
  wire \picorv32_core/n170 ;
  wire \picorv32_core/n180 ;
  wire \picorv32_core/n25 ;
  wire \picorv32_core/n274 ;
  wire \picorv32_core/n289_lutinv ;
  wire \picorv32_core/n304_lutinv ;
  wire \picorv32_core/n308_lutinv ;
  wire \picorv32_core/n328_lutinv ;
  wire \picorv32_core/n345 ;
  wire \picorv32_core/n407 ;
  wire \picorv32_core/n447 ;
  wire \picorv32_core/n456_0_al_n603 ;
  wire \picorv32_core/n456_1_al_n604 ;
  wire \picorv32_core/n472 ;
  wire \picorv32_core/n523_lutinv ;
  wire \picorv32_core/n524$4$_en ;
  wire \picorv32_core/n524$4$_en_al_n602 ;
  wire \picorv32_core/n554 ;
  wire \picorv32_core/n580 ;
  wire \picorv32_core/n662 ;
  wire \picorv32_core/n663 ;
  wire \picorv32_core/n664_lutinv ;
  wire \picorv32_core/n664_lutinv_placeOpt_1 ;
  wire \picorv32_core/n664_lutinv_placeOpt_2 ;
  wire \picorv32_core/n664_lutinv_placeOpt_3 ;
  wire \picorv32_core/n664_lutinv_placeOpt_4 ;
  wire \picorv32_core/n664_lutinv_placeOpt_5 ;
  wire \picorv32_core/n664_lutinv_placeOpt_6 ;
  wire \picorv32_core/n664_lutinv_placeOpt_7 ;
  wire \picorv32_core/n665_lutinv ;
  wire \picorv32_core/n666_lutinv ;
  wire \picorv32_core/n667_lutinv ;
  wire \picorv32_core/n668_lutinv ;
  wire \picorv32_core/n669_lutinv ;
  wire \picorv32_core/n669_lutinv_placeOpt_1 ;
  wire \picorv32_core/n669_lutinv_placeOpt_2 ;
  wire \picorv32_core/n669_lutinv_placeOpt_3 ;
  wire \picorv32_core/n669_lutinv_placeOpt_4 ;
  wire \picorv32_core/n728 ;
  wire \picorv32_core/n729 ;
  wire \picorv32_core/n731 ;
  wire \picorv32_core/n734_lutinv ;
  wire \picorv32_core/n746_lutinv ;
  wire \picorv32_core/n747 ;
  wire \picorv32_core/n98_lutinv ;
  wire \picorv32_core/pcpi_rs1$0$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$1$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$10$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$11$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$12$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$13$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$14$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$15$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$16$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$17$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$18$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$19$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$2$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$20$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$21$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$22$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$23$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$24$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$25$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$26$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$27$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$28$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$29$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$3$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$30$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$31$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$4$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$5$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$6$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$7$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$8$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$9$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs2$10$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$11$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$12$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$13$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$14$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$15$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$16$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$17$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$18$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$19$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$20$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$21$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$22$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$23$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$24$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$25$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$26$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$27$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$28$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$29$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$30$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$31$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$8$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$9$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/prefetched_high_word ;  // ../src/picorv32.v(329)
  wire \picorv32_core/sel15_b0_sel_is_3_o ;
  wire \picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ;
  wire \picorv32_core/sel15_b0_sel_is_3_o_placeOpt_2 ;
  wire \picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 ;
  wire \picorv32_core/sel39_b0_sel_is_3_o ;
  wire \picorv32_core/sel40_b0/or_or_B4_B5_o_or_B6__o_lutinv ;
  wire \picorv32_core/sel40_b1/or_or_B4_B5_o_or_B6__o_lutinv ;
  wire \picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv ;
  wire \picorv32_core/sub0/c1 ;
  wire \picorv32_core/sub0/c11 ;
  wire \picorv32_core/sub0/c13 ;
  wire \picorv32_core/sub0/c15 ;
  wire \picorv32_core/sub0/c17 ;
  wire \picorv32_core/sub0/c19 ;
  wire \picorv32_core/sub0/c21 ;
  wire \picorv32_core/sub0/c23 ;
  wire \picorv32_core/sub0/c25 ;
  wire \picorv32_core/sub0/c27 ;
  wire \picorv32_core/sub0/c29 ;
  wire \picorv32_core/sub0/c3 ;
  wire \picorv32_core/sub0/c31 ;
  wire \picorv32_core/sub0/c5 ;
  wire \picorv32_core/sub0/c7 ;
  wire \picorv32_core/sub0/c9 ;
  wire \picorv32_core/sub1/c1 ;
  wire \picorv32_core/sub1/c3 ;
  wire \picorv32_core/sub2/c1 ;
  wire \picorv32_core/sub2/c3 ;
  wire \picorv32_core/u179_sel_is_0_o ;
  wire \picorv32_core/u449_sel_is_0_o ;
  wire \picorv32_core/u616_sel_is_2_o ;
  wire \picorv32_core/u617_sel_is_2_o ;
  wire \picorv32_core/u625_sel_is_2_o ;
  wire resetn;  // ../src/top.v(33)
  wire resetn_i_pad;  // ../src/top.v(5)
  wire resetn_placeOpt_1;
  wire resetn_placeOpt_10;
  wire resetn_placeOpt_11;
  wire resetn_placeOpt_12;
  wire resetn_placeOpt_13;
  wire resetn_placeOpt_14;
  wire resetn_placeOpt_15;
  wire resetn_placeOpt_16;
  wire resetn_placeOpt_17;
  wire resetn_placeOpt_2;
  wire resetn_placeOpt_3;
  wire resetn_placeOpt_4;
  wire resetn_placeOpt_5;
  wire resetn_placeOpt_6;
  wire resetn_placeOpt_7;
  wire resetn_placeOpt_8;
  wire resetn_placeOpt_9;
  wire rxd_pad;  // ../src/top.v(14)
  wire trap_pad;  // ../src/top.v(6)
  wire txd_pad;  // ../src/top.v(13)
  wire \uart/add0/c1 ;
  wire \uart/add0/c11 ;
  wire \uart/add0/c13 ;
  wire \uart/add0/c15 ;
  wire \uart/add0/c17 ;
  wire \uart/add0/c19 ;
  wire \uart/add0/c21 ;
  wire \uart/add0/c23 ;
  wire \uart/add0/c25 ;
  wire \uart/add0/c27 ;
  wire \uart/add0/c29 ;
  wire \uart/add0/c3 ;
  wire \uart/add0/c31 ;
  wire \uart/add0/c5 ;
  wire \uart/add0/c7 ;
  wire \uart/add0/c9 ;
  wire \uart/add1/c1 ;
  wire \uart/add1/c3 ;
  wire \uart/add2/c1 ;
  wire \uart/add2/c3 ;
  wire \uart/add3/c1 ;
  wire \uart/add3/c3 ;
  wire \uart/lt0_c1 ;
  wire \uart/lt0_c11 ;
  wire \uart/lt0_c13 ;
  wire \uart/lt0_c15 ;
  wire \uart/lt0_c17 ;
  wire \uart/lt0_c19 ;
  wire \uart/lt0_c21 ;
  wire \uart/lt0_c23 ;
  wire \uart/lt0_c25 ;
  wire \uart/lt0_c27 ;
  wire \uart/lt0_c29 ;
  wire \uart/lt0_c3 ;
  wire \uart/lt0_c31 ;
  wire \uart/lt0_c5 ;
  wire \uart/lt0_c7 ;
  wire \uart/lt0_c9 ;
  wire \uart/mux12_b0_sel_is_3_o ;
  wire \uart/mux14_b0_sel_is_1_o ;
  wire \uart/mux15_b0_sel_is_2_o ;
  wire \uart/mux37_b0_sel_is_3_o ;
  wire \uart/mux51_b0_sel_is_3_o ;
  wire \uart/mux9_b0_sel_is_3_o ;
  wire \uart/n2 ;
  wire \uart/n30 ;
  wire \uart/n51_lutinv ;
  wire \uart/n9_lutinv ;
  wire \uart/sub1/c1 ;
  wire \uart/sub1/c3 ;
  wire \uart/u7_sel_is_3_o ;
  wire \uart/uart_op_clock ;  // ../src/uart.v(34)
  wire \uart/uart_status_fe ;  // ../src/uart.v(39)
  wire \uart/uart_status_rx ;  // ../src/uart.v(40)
  wire \uart/uart_status_rx_clr ;  // ../src/uart.v(156)
  wire \uart/uart_trigger_tx ;  // ../src/uart.v(44)
  wire uart_sel_lutinv;  // ../src/top.v(97)
  wire uart_sel_lutinv_placeOpt_1;
  wire uart_sel_lutinv_placeOpt_2;
  wire uart_sel_lutinv_placeOpt_3;

  EG_PHY_MSLICE #(
    //.LUT0("(~C*B)"),
    //.LUT1("(B*~D)"),
    .INIT_LUT0(16'b0000110000001100),
    .INIT_LUT1(16'b0000000011001100),
    .MODE("LOGIC"))
    \_al_u1000|_al_u1062  (
    .b({\picorv32_core/n663 ,\picorv32_core/n663 }),
    .c({open_n2,_al_u1061_o}),
    .d({_al_u999_o,open_n5}),
    .f({\picorv32_core/cpuregs_wrdata [9],\picorv32_core/cpuregs_wrdata [0]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("0"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1002|_al_u1001  (
    .a({open_n24,\picorv32_core/n450 [8]}),
    .b({open_n25,\picorv32_core/latched_branch }),
    .c({open_n26,\picorv32_core/latched_stalu }),
    .d({_al_u1001_o,\picorv32_core/reg_out [8]}),
    .e({\picorv32_core/n663 ,\picorv32_core/alu_out_q [8]}),
    .f({\picorv32_core/cpuregs_wrdata [8],_al_u1001_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+~A*B*~C*D+~A*B*C*D"),
    //.LUTG0("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011110000),
    .INIT_LUTF1(16'b0100010001110111),
    .INIT_LUTG0(16'b1111110011111010),
    .INIT_LUTG1(16'b0100011101000111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1003|picorv32_core/reg14_b7  (
    .a({\picorv32_core/n450 [7],\picorv32_core/n434 [7]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/n433 [7]}),
    .c({\picorv32_core/alu_out_q [7],_al_u885_o}),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [7],\picorv32_core/instr_sub }),
    .e({\picorv32_core/latched_stalu ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u1003_o,open_n65}),
    .q({open_n69,\picorv32_core/alu_out_q [7]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~C)"),
    //.LUT1("(B*~A)"),
    .INIT_LUT0(16'b0000110000001100),
    .INIT_LUT1(16'b0100010001000100),
    .MODE("LOGIC"))
    \_al_u1004|_al_u1060  (
    .a({_al_u1003_o,open_n70}),
    .b({\picorv32_core/n663 ,\picorv32_core/n663 }),
    .c({open_n71,_al_u1059_o}),
    .f({\picorv32_core/cpuregs_wrdata [7],\picorv32_core/cpuregs_wrdata [1]}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+~A*B*~C*D+~A*B*C*D"),
    //.LUTG0("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011110000),
    .INIT_LUTF1(16'b0100010001110111),
    .INIT_LUTG0(16'b1111110011111010),
    .INIT_LUTG1(16'b0100011101000111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1005|picorv32_core/reg14_b6  (
    .a({\picorv32_core/n450 [6],\picorv32_core/n434 [6]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/n433 [6]}),
    .c({\picorv32_core/alu_out_q [6],_al_u883_o}),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [6],\picorv32_core/instr_sub }),
    .e({\picorv32_core/latched_stalu ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u1005_o,open_n110}),
    .q({open_n114,\picorv32_core/alu_out_q [6]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~B)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0011000000110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0011000000110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1006|_al_u1054  (
    .b({open_n117,_al_u1053_o}),
    .c({\picorv32_core/n663 ,\picorv32_core/n663 }),
    .d({_al_u1005_o,open_n120}),
    .f({\picorv32_core/cpuregs_wrdata [6],\picorv32_core/cpuregs_wrdata [12]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("0"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1008|_al_u1007  (
    .a({_al_u1007_o,\picorv32_core/n450 [5]}),
    .b({open_n143,\picorv32_core/latched_branch }),
    .c({open_n144,\picorv32_core/latched_stalu }),
    .d({open_n147,\picorv32_core/reg_out [5]}),
    .e({\picorv32_core/n663 ,\picorv32_core/alu_out_q [5]}),
    .f({\picorv32_core/cpuregs_wrdata [5],_al_u1007_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1009 (
    .a({\picorv32_core/n450 [4],\picorv32_core/n450 [4]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [4],\picorv32_core/reg_out [4]}),
    .mi({open_n180,\picorv32_core/alu_out_q [4]}),
    .fx({open_n185,_al_u1009_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000111100001111),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1010|_al_u1052  (
    .a({_al_u1009_o,open_n188}),
    .c({open_n191,_al_u1051_o}),
    .e({\picorv32_core/n663 ,\picorv32_core/n663 }),
    .f({\picorv32_core/cpuregs_wrdata [4],\picorv32_core/cpuregs_wrdata [13]}));
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1011 (
    .a({\picorv32_core/n450 [31],\picorv32_core/n450 [31]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [31],\picorv32_core/reg_out [31]}),
    .mi({open_n228,\picorv32_core/alu_out_q [31]}),
    .fx({open_n233,_al_u1011_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~C)"),
    //.LUT1("(A*~D)"),
    .INIT_LUT0(16'b0000101000001010),
    .INIT_LUT1(16'b0000000010101010),
    .MODE("LOGIC"))
    \_al_u1012|_al_u1046  (
    .a({\picorv32_core/n663 ,\picorv32_core/n663 }),
    .c({open_n238,_al_u1045_o}),
    .d({_al_u1011_o,open_n241}),
    .f({\picorv32_core/cpuregs_wrdata [31],\picorv32_core/cpuregs_wrdata [16]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("(B*~D)"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("(B*~D)"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0000000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1014|_al_u1013  (
    .a({open_n260,\picorv32_core/n450 [30]}),
    .b({\picorv32_core/n663 ,\picorv32_core/latched_branch }),
    .c({open_n261,\picorv32_core/latched_stalu }),
    .d({_al_u1013_o,\picorv32_core/reg_out [30]}),
    .e({open_n264,\picorv32_core/alu_out_q [30]}),
    .f({\picorv32_core/cpuregs_wrdata [30],_al_u1013_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("0"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1016|_al_u1015  (
    .a({open_n285,\picorv32_core/n450 [3]}),
    .b({open_n286,\picorv32_core/latched_branch }),
    .c({open_n287,\picorv32_core/latched_stalu }),
    .d({_al_u1015_o,\picorv32_core/reg_out [3]}),
    .e({\picorv32_core/n663 ,\picorv32_core/alu_out_q [3]}),
    .f({\picorv32_core/cpuregs_wrdata [3],_al_u1015_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1017 (
    .a({\picorv32_core/n450 [29],\picorv32_core/n450 [29]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [29],\picorv32_core/reg_out [29]}),
    .mi({open_n322,\picorv32_core/alu_out_q [29]}),
    .fx({open_n327,_al_u1017_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~C)"),
    //.LUT1("(A*~C)"),
    .INIT_LUT0(16'b0000101000001010),
    .INIT_LUT1(16'b0000101000001010),
    .MODE("LOGIC"))
    \_al_u1018|_al_u1044  (
    .a({\picorv32_core/n663 ,\picorv32_core/n663 }),
    .c({_al_u1017_o,_al_u1043_o}),
    .f({\picorv32_core/cpuregs_wrdata [29],\picorv32_core/cpuregs_wrdata [17]}));
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1019 (
    .a({\picorv32_core/n450 [28],\picorv32_core/n450 [28]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [28],\picorv32_core/reg_out [28]}),
    .mi({open_n366,\picorv32_core/alu_out_q [28]}),
    .fx({open_n371,_al_u1019_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000011111111),
    .INIT_LUTG1(16'b0011001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1020|_al_u1038  (
    .b({_al_u1019_o,open_n376}),
    .d({open_n381,_al_u1037_o}),
    .e({\picorv32_core/n663 ,\picorv32_core/n663 }),
    .f({\picorv32_core/cpuregs_wrdata [28],\picorv32_core/cpuregs_wrdata [2]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("0"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1022|_al_u1021  (
    .a({_al_u1021_o,\picorv32_core/n450 [27]}),
    .b({open_n402,\picorv32_core/latched_branch }),
    .c({open_n403,\picorv32_core/latched_stalu }),
    .d({open_n406,\picorv32_core/reg_out [27]}),
    .e({\picorv32_core/n663 ,\picorv32_core/alu_out_q [27]}),
    .f({\picorv32_core/cpuregs_wrdata [27],_al_u1021_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("(A*~D)"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("(A*~D)"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0000000010101010),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1024|_al_u1023  (
    .a({\picorv32_core/n663 ,\picorv32_core/n450 [26]}),
    .b({open_n427,\picorv32_core/latched_branch }),
    .c({open_n428,\picorv32_core/latched_stalu }),
    .d({_al_u1023_o,\picorv32_core/reg_out [26]}),
    .e({open_n431,\picorv32_core/alu_out_q [26]}),
    .f({\picorv32_core/cpuregs_wrdata [26],_al_u1023_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1025 (
    .a({\picorv32_core/n450 [25],\picorv32_core/n450 [25]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [25],\picorv32_core/reg_out [25]}),
    .mi({open_n464,\picorv32_core/alu_out_q [25]}),
    .fx({open_n469,_al_u1025_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("0"),
    //.LUTG0("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0101010101010101),
    .INIT_LUTG1(16'b0011001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1026|_al_u1036  (
    .a({open_n472,_al_u1035_o}),
    .b({_al_u1025_o,open_n473}),
    .e({\picorv32_core/n663 ,\picorv32_core/n663 }),
    .f({\picorv32_core/cpuregs_wrdata [25],\picorv32_core/cpuregs_wrdata [20]}));
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1027 (
    .a({\picorv32_core/n450 [24],\picorv32_core/n450 [24]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [24],\picorv32_core/reg_out [24]}),
    .mi({open_n512,\picorv32_core/alu_out_q [24]}),
    .fx({open_n517,_al_u1027_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~D)"),
    //.LUT1("(B*~D)"),
    .INIT_LUT0(16'b0000000011001100),
    .INIT_LUT1(16'b0000000011001100),
    .MODE("LOGIC"))
    \_al_u1028|_al_u1034  (
    .b({\picorv32_core/n663 ,\picorv32_core/n663 }),
    .d({_al_u1027_o,_al_u1033_o}),
    .f({\picorv32_core/cpuregs_wrdata [24],\picorv32_core/cpuregs_wrdata [21]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("0"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1030|_al_u1029  (
    .a({_al_u1029_o,\picorv32_core/n450 [23]}),
    .b({open_n544,\picorv32_core/latched_branch }),
    .c({open_n545,\picorv32_core/latched_stalu }),
    .d({open_n548,\picorv32_core/reg_out [23]}),
    .e({\picorv32_core/n663 ,\picorv32_core/alu_out_q [23]}),
    .f({\picorv32_core/cpuregs_wrdata [23],_al_u1029_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("(B*~A)"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("(B*~A)"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0100010001000100),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0100010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1032|_al_u1031  (
    .a({_al_u1031_o,\picorv32_core/n450 [22]}),
    .b({\picorv32_core/n663 ,\picorv32_core/latched_branch }),
    .c({open_n569,\picorv32_core/latched_stalu }),
    .d({open_n572,\picorv32_core/reg_out [22]}),
    .e({open_n573,\picorv32_core/alu_out_q [22]}),
    .f({\picorv32_core/cpuregs_wrdata [22],_al_u1031_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1033 (
    .a({\picorv32_core/n450 [21],\picorv32_core/n450 [21]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [21],\picorv32_core/reg_out [21]}),
    .mi({open_n606,\picorv32_core/alu_out_q [21]}),
    .fx({open_n611,_al_u1033_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1035 (
    .a({\picorv32_core/n450 [20],\picorv32_core/n450 [20]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [20],\picorv32_core/reg_out [20]}),
    .mi({open_n626,\picorv32_core/alu_out_q [20]}),
    .fx({open_n631,_al_u1035_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*B*C*D"),
    //.LUTG0("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+~A*B*~C*D+~A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011110000),
    .INIT_LUTF1(16'b0100011101000111),
    .INIT_LUTG0(16'b1111110011111010),
    .INIT_LUTG1(16'b0100010001110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1037|picorv32_core/reg14_b2  (
    .a({\picorv32_core/n450 [2],\picorv32_core/n434 [2]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/n433 [2]}),
    .c({\picorv32_core/reg_out [2],_al_u851_o}),
    .clk(clk_pad),
    .d({\picorv32_core/alu_out_q [2],\picorv32_core/instr_sub }),
    .e({\picorv32_core/latched_stalu ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u1037_o,open_n650}),
    .q({open_n654,\picorv32_core/alu_out_q [2]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("(B*~A)"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("(B*~A)"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0100010001000100),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0100010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1040|_al_u1039  (
    .a({_al_u1039_o,\picorv32_core/n450 [19]}),
    .b({\picorv32_core/n663 ,\picorv32_core/latched_branch }),
    .c({open_n655,\picorv32_core/latched_stalu }),
    .d({open_n658,\picorv32_core/reg_out [19]}),
    .e({open_n659,\picorv32_core/alu_out_q [19]}),
    .f({\picorv32_core/cpuregs_wrdata [19],_al_u1039_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("(B*~D)"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("(B*~D)"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0000000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1042|_al_u1041  (
    .a({open_n680,\picorv32_core/n450 [18]}),
    .b({\picorv32_core/n663 ,\picorv32_core/latched_branch }),
    .c({open_n681,\picorv32_core/latched_stalu }),
    .d({_al_u1041_o,\picorv32_core/reg_out [18]}),
    .e({open_n684,\picorv32_core/alu_out_q [18]}),
    .f({\picorv32_core/cpuregs_wrdata [18],_al_u1041_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1043 (
    .a({\picorv32_core/n450 [17],\picorv32_core/n450 [17]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [17],\picorv32_core/reg_out [17]}),
    .mi({open_n717,\picorv32_core/alu_out_q [17]}),
    .fx({open_n722,_al_u1043_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1045 (
    .a({\picorv32_core/n450 [16],\picorv32_core/n450 [16]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [16],\picorv32_core/reg_out [16]}),
    .mi({open_n737,\picorv32_core/alu_out_q [16]}),
    .fx({open_n742,_al_u1045_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("(B*~A)"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("(B*~A)"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0100010001000100),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0100010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1048|_al_u1047  (
    .a({_al_u1047_o,\picorv32_core/n450 [15]}),
    .b({\picorv32_core/n663 ,\picorv32_core/latched_branch }),
    .c({open_n745,\picorv32_core/latched_stalu }),
    .d({open_n748,\picorv32_core/reg_out [15]}),
    .e({open_n749,\picorv32_core/alu_out_q [15]}),
    .f({\picorv32_core/cpuregs_wrdata [15],_al_u1047_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("(D*~A)"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("(D*~A)"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0101010100000000),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0101010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1050|_al_u1049  (
    .a({_al_u1049_o,\picorv32_core/n450 [14]}),
    .b({open_n770,\picorv32_core/latched_branch }),
    .c({open_n771,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/n663 ,\picorv32_core/reg_out [14]}),
    .e({open_n774,\picorv32_core/alu_out_q [14]}),
    .f({\picorv32_core/cpuregs_wrdata [14],_al_u1049_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1051 (
    .a({\picorv32_core/n450 [13],\picorv32_core/n450 [13]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [13],\picorv32_core/reg_out [13]}),
    .mi({open_n807,\picorv32_core/alu_out_q [13]}),
    .fx({open_n812,_al_u1051_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1053 (
    .a({\picorv32_core/n450 [12],\picorv32_core/n450 [12]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [12],\picorv32_core/reg_out [12]}),
    .mi({open_n827,\picorv32_core/alu_out_q [12]}),
    .fx({open_n832,_al_u1053_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("0"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1056|_al_u1055  (
    .a({_al_u1055_o,\picorv32_core/n450 [11]}),
    .b({open_n835,\picorv32_core/latched_branch }),
    .c({open_n836,\picorv32_core/latched_stalu }),
    .d({open_n839,\picorv32_core/reg_out [11]}),
    .e({\picorv32_core/n663 ,\picorv32_core/alu_out_q [11]}),
    .f({\picorv32_core/cpuregs_wrdata [11],_al_u1055_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUTF1("(B*~D)"),
    //.LUTG0("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    //.LUTG1("(B*~D)"),
    .INIT_LUTF0(16'b0111010001110111),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b0100010001000111),
    .INIT_LUTG1(16'b0000000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1058|_al_u1057  (
    .a({open_n860,\picorv32_core/n450 [10]}),
    .b({\picorv32_core/n663 ,\picorv32_core/latched_branch }),
    .c({open_n861,\picorv32_core/latched_stalu }),
    .d({_al_u1057_o,\picorv32_core/reg_out [10]}),
    .e({open_n864,\picorv32_core/alu_out_q [10]}),
    .f({\picorv32_core/cpuregs_wrdata [10],_al_u1057_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+~A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011110000),
    .INIT_LUTF1(16'b1101110011011111),
    .INIT_LUTG0(16'b1111110011111010),
    .INIT_LUTG1(16'b0001000000010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1059|picorv32_core/reg14_b1  (
    .a({\picorv32_core/alu_out_q [1],\picorv32_core/n434 [1]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/n433 [1]}),
    .c({\picorv32_core/latched_stalu ,_al_u829_o}),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [1],\picorv32_core/instr_sub }),
    .e({\picorv32_core/n450 [1],\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u1059_o,open_n901}),
    .q({open_n905,\picorv32_core/alu_out_q [1]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1061 (
    .a({\picorv32_core/n450 [0],\picorv32_core/n450 [0]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [0],\picorv32_core/reg_out [0]}),
    .mi({open_n918,\picorv32_core/alu_out_q [0]}),
    .fx({open_n923,_al_u1061_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(0*D*~C*B*~A)"),
    //.LUT1("(1*B*~A*D*~C)"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000010000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1063 (
    .a({\uart/uart_status_rxd [2],\uart/uart_status_rxd [0]}),
    .b({\uart/uart_status_rxd [3],\uart/uart_status_rxd [1]}),
    .c({\uart/uart_status_rxd [0],\uart/uart_status_rxd [2]}),
    .d({\uart/uart_status_rxd [1],\uart/uart_status_rxd [3]}),
    .mi({open_n938,\uart/uart_op_clock }),
    .fx({open_n943,_al_u1063_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~D*~(0*~(~C*B)))"),
    //.LUTF1("0"),
    //.LUTG0("(~A*~D*~(1*~(~C*B)))"),
    //.LUTG1("D*A*~B*~C+D*A*B*~C"),
    .INIT_LUTF0(16'b0000000001010101),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000100),
    .INIT_LUTG1(16'b0000101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1066|_al_u1067  (
    .a({rxd_pad,\uart/uart_status_rxd [3]}),
    .b({open_n946,_al_u1065_o}),
    .c({\uart/uart_status_rxd [0],\uart/uart_status_rxd [0]}),
    .d({_al_u1065_o,_al_u1066_o}),
    .e(\uart/uart_cnt_rx [2:1]),
    .f({_al_u1066_o,_al_u1067_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*~D))"),
    //.LUTF1("0"),
    //.LUTG0("(~B*~(~C*~D))"),
    //.LUTG1("C*~D*~B*~A+C*~D*~B*A"),
    .INIT_LUTF0(16'b0011001100110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0011001100110000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1071|_al_u1165  (
    .b({\uart/uart_cnt_rx [1],\uart/uart_status_rxd [3]}),
    .c({rxd_pad,rxd_pad}),
    .d({\uart/uart_status_rxd [0],\uart/uart_status_rxd [0]}),
    .e({_al_u1070_o,open_n973}),
    .f({_al_u1071_o,_al_u1165_o}));
  // ../src/uart.v(263)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~((B*~(D)*~(0)+~(B)*D*~(0)+~(B)*D*0))*~(C)+~A*(B*~(D)*~(0)+~(B)*D*~(0)+~(B)*D*0)*~(C)+~(~A)*(B*~(D)*~(0)+~(B)*D*~(0)+~(B)*D*0)*C+~A*(B*~(D)*~(0)+~(B)*D*~(0)+~(B)*D*0)*C)"),
    //.LUTF1("~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D"),
    //.LUTG0("(~A*~((B*~(D)*~(1)+~(B)*D*~(1)+~(B)*D*1))*~(C)+~A*(B*~(D)*~(1)+~(B)*D*~(1)+~(B)*D*1)*~(C)+~(~A)*(B*~(D)*~(1)+~(B)*D*~(1)+~(B)*D*1)*C+~A*(B*~(D)*~(1)+~(B)*D*~(1)+~(B)*D*1)*C)"),
    //.LUTG1("~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011010111000101),
    .INIT_LUTF1(16'b0111111101111100),
    .INIT_LUTG0(16'b0011010100000101),
    .INIT_LUTG1(16'b1111111111001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1074|uart/reg8_b0  (
    .a({rxd_pad,_al_u1074_o}),
    .b({\uart/uart_cnt_rx [0],_al_u1068_o}),
    .c({_al_u1065_o,\uart/uart_status_rxd [3]}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d(\uart/uart_cnt_rx [1:0]),
    .e({\uart/uart_status_rxd [0],\uart/uart_cnt_rx [1]}),
    .sr(resetn_placeOpt_9),
    .f({_al_u1074_o,open_n1008}),
    .q({open_n1012,\uart/uart_cnt_rx [0]}));  // ../src/uart.v(263)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+~(A)*B*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+A*~(B)*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+A*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0+A*B*C*D*0)"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+~(A)*B*~(C)*~(D)*~(1)+A*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+A*~(B)*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+A*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+A*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1+A*B*C*D*1)"),
    //.LUTG1("A*~B*~C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b1010111110100111),
    .INIT_LUTF1(16'b0010111011001100),
    .INIT_LUTG0(16'b1111111111101111),
    .INIT_LUTG1(16'b0010001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1077|_al_u1081  (
    .a({_al_u1076_o,_al_u1076_o}),
    .b({\uart/uart_status_txd [3],\uart/uart_status_txd [0]}),
    .c({\uart/uart_status_txd [0],\uart/uart_status_txd [1]}),
    .d({\uart/uart_status_txd [1],\uart/uart_status_txd [2]}),
    .e({\uart/uart_status_txd [2],\uart/uart_status_txd [3]}),
    .f({_al_u1077_o,_al_u1081_o}));
  // ../src/uart.v(145)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~C*D*~B+A*C*D*~B+~A*~C*~D*B+A*~C*~D*B+~A*C*~D*B+A*C*~D*B+A*~C*D*B+A*C*D*B"),
    //.LUTF1("(A@(~D*~B))"),
    //.LUTG0("0"),
    //.LUTG1("(A@(~D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011001100),
    .INIT_LUTF1(16'b1010101010011001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1010101010011001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1079|uart/reg4_b2  (
    .a({\uart/uart_status_txd [3],\uart/n35 [2]}),
    .b({\uart/uart_status_txd [1],\uart/uart_status_txd [2]}),
    .ce(\uart/n30 ),
    .clk(clk_pad),
    .d({\uart/uart_status_txd [2],_al_u1076_o}),
    .e({open_n1037,_al_u1079_o}),
    .sr(resetn_placeOpt_1),
    .f({_al_u1079_o,open_n1052}),
    .q({open_n1056,\uart/uart_status_txd [2]}));  // ../src/uart.v(145)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~D)"),
    //.LUT1("(C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011111111),
    .INIT_LUT1(16'b0010000000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1084|picorv32_core/mem_do_prefetch_reg  (
    .a({\picorv32_core/sel39_b0_sel_is_3_o ,open_n1057}),
    .b({\picorv32_core/instr_jal ,open_n1058}),
    .c({resetn_placeOpt_11,open_n1059}),
    .ce(\picorv32_core/u617_sel_is_2_o ),
    .clk(clk_pad),
    .d({open_n1060,\picorv32_core/instr_jalr }),
    .sr(\picorv32_core/n747 ),
    .f({\picorv32_core/u617_sel_is_2_o ,open_n1073}),
    .q({open_n1077,\picorv32_core/mem_do_prefetch }));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~B)"),
    //.LUT1("(D*~A*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001100110011),
    .INIT_LUT1(16'b0101000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1084|picorv32_core/mem_do_prefetch_reg_placeOpt_1  (
    .a({\picorv32_core/instr_jal ,open_n1078}),
    .b({open_n1079,\picorv32_core/instr_jalr }),
    .c({\picorv32_core/sel39_b0_sel_is_3_o ,open_n1080}),
    .ce(\picorv32_core/u617_sel_is_2_o ),
    .clk(clk_pad),
    .d({resetn_placeOpt_11,open_n1081}),
    .sr(\picorv32_core/n747 ),
    .q({open_n1099,\picorv32_core/mem_do_prefetch_placeOpt_1 }));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~B)"),
    //.LUT1("(C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001100110011),
    .INIT_LUT1(16'b0010000000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1084|picorv32_core/mem_do_prefetch_reg_placeOpt_2  (
    .a({\picorv32_core/sel39_b0_sel_is_3_o ,open_n1100}),
    .b({\picorv32_core/instr_jal ,\picorv32_core/instr_jalr }),
    .c({resetn_placeOpt_11,open_n1101}),
    .ce(\picorv32_core/u617_sel_is_2_o ),
    .clk(clk_pad),
    .sr(\picorv32_core/n747 ),
    .q({open_n1121,\picorv32_core/mem_do_prefetch_placeOpt_2 }));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~C)"),
    //.LUT1("(A*~B*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100001111),
    .INIT_LUT1(16'b0010000000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1084|picorv32_core/mem_do_prefetch_reg_placeOpt_3  (
    .a({resetn_placeOpt_11,open_n1122}),
    .b({\picorv32_core/instr_jal ,open_n1123}),
    .c({\picorv32_core/sel39_b0_sel_is_3_o ,\picorv32_core/instr_jalr }),
    .ce(\picorv32_core/u617_sel_is_2_o ),
    .clk(clk_pad),
    .sr(\picorv32_core/n747 ),
    .q({open_n1143,\picorv32_core/mem_do_prefetch_placeOpt_3 }));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~B)"),
    //.LUT1("(A*~D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001100110011),
    .INIT_LUT1(16'b0000000010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1084|picorv32_core/mem_do_prefetch_reg_placeOpt_4  (
    .a({resetn_placeOpt_11,open_n1144}),
    .b({open_n1145,\picorv32_core/instr_jalr }),
    .c({\picorv32_core/sel39_b0_sel_is_3_o ,open_n1146}),
    .ce(\picorv32_core/u617_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_jal ,open_n1147}),
    .sr(\picorv32_core/n747 ),
    .q({open_n1165,\picorv32_core/mem_do_prefetch_placeOpt_4 }));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~D)"),
    //.LUT1("(A*~B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011111111),
    .INIT_LUT1(16'b0010001000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1084|picorv32_core/mem_do_prefetch_reg_placeOpt_5  (
    .a({resetn_placeOpt_11,open_n1166}),
    .b({\picorv32_core/instr_jal ,open_n1167}),
    .ce(\picorv32_core/u617_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/sel39_b0_sel_is_3_o ,\picorv32_core/instr_jalr }),
    .sr(\picorv32_core/n747 ),
    .q({open_n1187,\picorv32_core/mem_do_prefetch_placeOpt_5 }));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~D)"),
    //.LUT1("(A*~B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011111111),
    .INIT_LUT1(16'b0010001000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1084|picorv32_core/mem_do_prefetch_reg_placeOpt_6  (
    .a({resetn_placeOpt_11,open_n1188}),
    .b({\picorv32_core/instr_jal ,open_n1189}),
    .ce(\picorv32_core/u617_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/sel39_b0_sel_is_3_o ,\picorv32_core/instr_jalr }),
    .sr(\picorv32_core/n747 ),
    .q({open_n1209,\picorv32_core/mem_do_prefetch_placeOpt_6 }));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~B)"),
    //.LUT1("(A*~D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001100110011),
    .INIT_LUT1(16'b0000000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1084|picorv32_core/mem_do_prefetch_reg_placeOpt_7  (
    .a({resetn_placeOpt_11,open_n1210}),
    .b({\picorv32_core/sel39_b0_sel_is_3_o ,\picorv32_core/instr_jalr }),
    .ce(\picorv32_core/u617_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_jal ,open_n1213}),
    .sr(\picorv32_core/n747 ),
    .q({open_n1231,\picorv32_core/mem_do_prefetch_placeOpt_7 }));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~C)"),
    //.LUT1("(C*~B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100001111),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1084|picorv32_core/mem_do_prefetch_reg_placeOpt_8  (
    .b({\picorv32_core/instr_jal ,open_n1234}),
    .c({resetn_placeOpt_11,\picorv32_core/instr_jalr }),
    .ce(\picorv32_core/u617_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/sel39_b0_sel_is_3_o ,open_n1235}),
    .sr(\picorv32_core/n747 ),
    .q({open_n1253,\picorv32_core/mem_do_prefetch_placeOpt_8 }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(~D*~A))"),
    //.LUT1("(~C*~B*~D)"),
    .INIT_LUT0(16'b0011111100101010),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"))
    \_al_u1086|_al_u1227  (
    .a({open_n1254,_al_u1068_o}),
    .b({\uart/uart_smp_rx [2],\uart/n51_lutinv }),
    .c({\uart/uart_smp_rx [3],_al_u1065_o}),
    .d({\uart/uart_smp_rx [1],\uart/uart_smp_rx [1]}),
    .f({_al_u1086_o,_al_u1227_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("(~A*~D*(0*~(B)*~(C)+0*B*~(C)+~(0)*B*C+0*B*C))"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("(~A*~D*(1*~(B)*~(C)+1*B*~(C)+~(1)*B*C+1*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b0000000001000000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b0000000001000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1088|picorv32_core/reg17_b1  (
    .a({\picorv32_core/mem_la_secondword ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 }),
    .b({\picorv32_core/reg_out [1],\picorv32_core/latched_stalu }),
    .c({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 ,\picorv32_core/reg_out [1]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({_al_u700_o_placeOpt_2,\picorv32_core/alu_out_q [1]}),
    .e({\picorv32_core/reg_next_pc [1],\picorv32_core/reg_next_pc [1]}),
    .sr(resetn_placeOpt_10),
    .f({_al_u1088_o,\picorv32_core/n500 [1]}),
    .q({open_n1292,\picorv32_core/reg_pc [1]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1241)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B*~(C*A))"),
    //.LUT1("(B*~A*~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000010011),
    .INIT_LUT1(16'b0000010000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1089|picorv32_core/clear_prefetched_high_word_q_reg  (
    .a({\picorv32_core/clear_prefetched_high_word_q ,\picorv32_core/clear_prefetched_high_word_q }),
    .b({\picorv32_core/prefetched_high_word ,\picorv32_core/n447 }),
    .c({\picorv32_core/n447 ,\picorv32_core/prefetched_high_word }),
    .ce(\picorv32_core/prefetched_high_word ),
    .clk(clk_pad),
    .d({_al_u1088_o,trap_pad}),
    .mi({open_n1303,1'b0}),
    .sr(\picorv32_core/n447 ),
    .f({_al_u1089_o,\picorv32_core/u179_sel_is_0_o }),
    .q({open_n1307,\picorv32_core/clear_prefetched_high_word_q }));  // ../src/picorv32.v(1241)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("~(~B*~(A*C))"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b1110110011101100),
    .MODE("LOGIC"))
    \_al_u1090|_al_u700  (
    .a({\picorv32_core/mem_do_rinst ,open_n1308}),
    .b({\picorv32_core/mem_valid ,\picorv32_core/mem_do_rinst }),
    .c({_al_u1089_o,open_n1309}),
    .d({open_n1312,\picorv32_core/mem_do_prefetch_placeOpt_1 }),
    .f({\picorv32_core/mem_xfer ,_al_u700_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~C)"),
    //.LUT1("~(~B*~(C*A))"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b1110110011101100),
    .MODE("LOGIC"))
    \_al_u1090|_al_u700_placeOpt_1  (
    .a({_al_u1089_o,\picorv32_core/mem_do_rinst }),
    .b({\picorv32_core/mem_valid ,open_n1331}),
    .c({\picorv32_core/mem_do_rinst ,\picorv32_core/mem_do_prefetch_placeOpt_1 }),
    .f({open_n1349,_al_u700_o_placeOpt_1}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A)"),
    //.LUT1("~(~D*~(C*A))"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b1111111110100000),
    .MODE("LOGIC"))
    \_al_u1090|_al_u700_placeOpt_1_al_u2582  (
    .a({_al_u1089_o,\picorv32_core/mem_do_prefetch_placeOpt_1 }),
    .c({\picorv32_core/mem_do_rinst ,\picorv32_core/mem_do_rinst }),
    .d({\picorv32_core/mem_valid ,open_n1359}),
    .f({\picorv32_core/mem_xfer_placeOpt_1 ,open_n1373}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("~(~C*~(A*D))"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b1111101011110000),
    .MODE("LOGIC"))
    \_al_u1090|_al_u700_placeOpt_2  (
    .a({\picorv32_core/mem_do_rinst ,\picorv32_core/mem_do_rinst }),
    .c({\picorv32_core/mem_valid ,open_n1381}),
    .d({_al_u1089_o,\picorv32_core/mem_do_prefetch_placeOpt_1 }),
    .f({open_n1397,_al_u700_o_placeOpt_2}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("~(~C*~(B*D))"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"))
    \_al_u1090|_al_u700_placeOpt_2_al_u2583  (
    .a({open_n1403,\picorv32_core/mem_do_prefetch_placeOpt_1 }),
    .b({\picorv32_core/mem_do_rinst ,\picorv32_core/mem_do_rinst }),
    .c({\picorv32_core/mem_valid ,open_n1404}),
    .d({_al_u1089_o,open_n1407}),
    .f({\picorv32_core/mem_xfer_placeOpt_2 ,open_n1421}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A)"),
    //.LUT1("~(~D*~(A*C))"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b1111111110100000),
    .MODE("LOGIC"))
    \_al_u1090|_al_u700_placeOpt_3  (
    .a({\picorv32_core/mem_do_rinst ,\picorv32_core/mem_do_prefetch_placeOpt_1 }),
    .c({_al_u1089_o,\picorv32_core/mem_do_rinst }),
    .d({\picorv32_core/mem_valid ,open_n1431}),
    .f({open_n1445,_al_u700_o_placeOpt_3}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("~(~A*~(B*D))"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b1110111010101010),
    .MODE("LOGIC"))
    \_al_u1090|_al_u700_placeOpt_3_al_u2584  (
    .a({\picorv32_core/mem_valid ,open_n1451}),
    .b({\picorv32_core/mem_do_rinst ,\picorv32_core/mem_do_rinst }),
    .d({_al_u1089_o,\picorv32_core/mem_do_prefetch_placeOpt_1 }),
    .f({\picorv32_core/mem_xfer_placeOpt_3 ,open_n1469}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("~(~C*~(B*A))"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b1111100011111000),
    .MODE("LOGIC"))
    \_al_u1090|_al_u700_placeOpt_4  (
    .a({_al_u1089_o,\picorv32_core/mem_do_rinst }),
    .b({\picorv32_core/mem_do_rinst ,\picorv32_core/mem_do_prefetch_placeOpt_1 }),
    .c({\picorv32_core/mem_valid ,open_n1475}),
    .f({\picorv32_core/mem_xfer_placeOpt_4 ,open_n1493}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~C)"),
    //.LUT1("~(~D*~(C*A))"),
    .INIT_LUT0(16'b0000001100000011),
    .INIT_LUT1(16'b1111111110100000),
    .MODE("LOGIC"))
    \_al_u1090|_al_u700_placeOpt_5  (
    .a({_al_u1089_o,open_n1499}),
    .b({open_n1500,\picorv32_core/mem_do_rinst }),
    .c({\picorv32_core/mem_do_rinst ,\picorv32_core/mem_do_prefetch_placeOpt_1 }),
    .d({\picorv32_core/mem_valid ,open_n1503}),
    .f({\picorv32_core/mem_xfer_placeOpt_5 ,open_n1517}));
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(C*A)"),
    //.LUT1("(~B*~D*~C*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010000010100000),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1091|picorv32_core/instr_slti_reg  (
    .a({\picorv32_core/n289_lutinv ,\picorv32_core/n289_lutinv }),
    .b({\picorv32_core/mem_rdata_q [19],open_n1523}),
    .c({\picorv32_core/mem_rdata_q [15],\picorv32_core/is_alu_reg_imm }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [16],open_n1524}),
    .sr(resetn_placeOpt_13),
    .f({_al_u1091_o,open_n1537}),
    .q({open_n1541,\picorv32_core/instr_slti }));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~A)"),
    //.LUTF1("0"),
    //.LUTG0("(~D*~A)"),
    //.LUTG1("~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000000001010101),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000001010101),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1094|_al_u1497  (
    .a({open_n1542,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({\picorv32_core/mem_rdata_q [4],open_n1543}),
    .c({\picorv32_core/mem_rdata_q [5],open_n1544}),
    .d({\picorv32_core/mem_rdata_q [6],\picorv32_core/mem_16bit_buffer [5]}),
    .e({_al_u1093_o,open_n1547}),
    .f({\picorv32_core/n328_lutinv ,_al_u1497_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*B*~C*~D+A*B*C*~D"),
    //.LUTF1("0"),
    //.LUTG0("0"),
    //.LUTG1("C*~B*~A*~D+C*B*~A*~D+C*~B*A*~D+C*B*A*~D+C*~B*~A*D+C*B*~A*D+C*~B*A*D+C*B*A*D"),
    .INIT_LUTF0(16'b0000000010001000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1095|_al_u1093  (
    .a({open_n1568,\picorv32_core/mem_rdata_q [0]}),
    .b({open_n1569,\picorv32_core/mem_rdata_q [1]}),
    .c({\picorv32_core/n328_lutinv ,open_n1570}),
    .d({open_n1573,\picorv32_core/mem_rdata_q [3]}),
    .e({_al_u1092_o,\picorv32_core/mem_rdata_q [2]}),
    .f({_al_u1095_o,_al_u1093_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~(D*~B))"),
    //.LUTF1("~D*~A*~C*~B+~D*~A*~C*B"),
    //.LUTG0("~(A*~(D*~B))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011101010101),
    .INIT_LUTF1(16'b0000000000000101),
    .INIT_LUTG0(16'b0111011101010101),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1096|picorv32_core/reg11_b3  (
    .a({\picorv32_core/mem_rdata_q [24],_al_u904_o}),
    .b({open_n1594,_al_u803_o}),
    .c({\picorv32_core/mem_rdata_q [22],open_n1595}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [23],\picorv32_core/mem_rdata_q [23]}),
    .e({\picorv32_core/mem_rdata_q [28],open_n1596}),
    .f({_al_u1096_o,open_n1612}),
    .q({open_n1616,\picorv32_core/decoded_imm [3]}));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~D*~A)"),
    //.LUTF1("0"),
    //.LUTG0("(~B*~D*~A)"),
    //.LUTG1("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+C*B*~A*~D"),
    .INIT_LUTF0(16'b0000000000010001),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000010001),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1097|_al_u973  (
    .a({\picorv32_core/mem_rdata_q [25],\picorv32_core/mem_rdata_q [25]}),
    .b({open_n1617,\picorv32_core/mem_rdata_q [27]}),
    .d({\picorv32_core/mem_rdata_q [26],\picorv32_core/mem_rdata_q [26]}),
    .e({_al_u1096_o,open_n1622}),
    .f({_al_u1097_o,_al_u973_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(0*D*~C*~B*A)"),
    //.LUT1("(1*B*~A*~D*C)"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000001000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1100 (
    .a({\picorv32_core/mem_rdata_q [29],_al_u1097_o}),
    .b({\picorv32_core/mem_rdata_q [30],\picorv32_core/mem_rdata_q [27]}),
    .c({_al_u1097_o,\picorv32_core/mem_rdata_q [29]}),
    .d({\picorv32_core/mem_rdata_q [27],\picorv32_core/mem_rdata_q [30]}),
    .mi({open_n1655,\picorv32_core/mem_rdata_q [31]}),
    .fx({open_n1660,_al_u1100_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(D*A)"),
    //.LUT1("(~A*~(~D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101000000000),
    .INIT_LUT1(16'b0101010100010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1102|picorv32_core/instr_srai_reg  (
    .a({\picorv32_core/n345 ,\picorv32_core/n345 }),
    .b({\picorv32_core/n304_lutinv ,open_n1663}),
    .c({\picorv32_core/mem_rdata_q [12],open_n1664}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [13],\picorv32_core/is_alu_reg_imm }),
    .f({_al_u1102_o,open_n1678}),
    .q({open_n1682,\picorv32_core/instr_srai }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(D*A)"),
    //.LUT1("(B*D*~(~C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101000000000),
    .INIT_LUT1(16'b1100100000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1105|picorv32_core/latched_compr_reg  (
    .a({\picorv32_core/latched_branch ,\picorv32_core/n663 }),
    .b({\picorv32_core/latched_rd [4],open_n1683}),
    .c({\picorv32_core/latched_store ,open_n1684}),
    .ce(\picorv32_core/u616_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/u616_sel_is_2_o ,resetn_placeOpt_7}),
    .mi({open_n1695,\picorv32_core/compressed_instr }),
    .f({\picorv32_core/n456_1_al_n604 ,\picorv32_core/u616_sel_is_2_o }),
    .q({open_n1700,\picorv32_core/latched_compr }));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*~A))"),
    //.LUT1("(~C*D*~(~A*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110001010000),
    .INIT_LUT1(16'b0000111000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1106|picorv32_core/reg24_b4  (
    .a({\picorv32_core/latched_store ,_al_u1153_o}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/n663 }),
    .c({\picorv32_core/latched_rd [4],\picorv32_core/latched_rd [4]}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/u616_sel_is_2_o ,\picorv32_core/decoded_rd [4]}),
    .f({\picorv32_core/n456_0_al_n603 ,open_n1714}),
    .q({open_n1718,\picorv32_core/latched_rd [4]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(~D*~B*~(~C*~A)))"),
    //.LUT1("(1*~(~D*~B*~(~C*~A)))"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1111111111001101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1107 (
    .a({\uart/uart_odr [6],\uart/uart_odr [6]}),
    .b({\uart/uart_status_txd [0],\uart/uart_status_txd [0]}),
    .c({\uart/uart_status_txd [1],\uart/uart_status_txd [1]}),
    .d({\uart/uart_status_txd [2],\uart/uart_status_txd [2]}),
    .mi({open_n1731,\uart/uart_status_txd [3]}),
    .fx({open_n1736,_al_u1107_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(~(B)*~(C)*~(D)*~(0)+~(B)*C*~(D)*~(0)+B*C*~(D)*~(0)+~(B)*~(C)*D*~(0)+B*~(C)*D*~(0)+~(B)*C*D*~(0)+B*C*D*~(0)+~(B)*~(C)*~(D)*0+~(B)*C*~(D)*0))"),
    //.LUT1("(A*(~(B)*~(C)*~(D)*~(1)+~(B)*C*~(D)*~(1)+B*C*~(D)*~(1)+~(B)*~(C)*D*~(1)+B*~(C)*D*~(1)+~(B)*C*D*~(1)+B*C*D*~(1)+~(B)*~(C)*~(D)*1+~(B)*C*~(D)*1))"),
    .INIT_LUT0(16'b1010101010100010),
    .INIT_LUT1(16'b0000000000100010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1108 (
    .a({_al_u1107_o,_al_u1107_o}),
    .b({\uart/uart_status_txd [0],\uart/uart_status_txd [0]}),
    .c({\uart/uart_status_txd [1],\uart/uart_status_txd [1]}),
    .d({\uart/uart_status_txd [2],\uart/uart_status_txd [2]}),
    .mi({open_n1751,txd_pad}),
    .fx({open_n1756,_al_u1108_o}));
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D)"),
    //.LUTF1("~A*~D*~B*~C+~A*D*~B*~C+~A*~D*B*~C+~A*D*B*~C+~A*~D*~B*C+~A*D*~B*C+~A*~D*B*C+~A*D*B*C"),
    //.LUTG0("(~D)"),
    //.LUTG1("~A*~D*~B*~C+~A*~D*B*~C+~A*D*B*~C+~A*~D*~B*C+~A*~D*B*C+~A*D*B*C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011111111),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000000011111111),
    .INIT_LUTG1(16'b0100010001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1109|uart/reg3_b7  (
    .a({_al_u1108_o,open_n1759}),
    .b({\uart/uart_odr [7],open_n1760}),
    .ce(\uart/mux15_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\uart/uart_status_txd [0],mem_la_wdata[7]}),
    .e({_al_u799_o,open_n1763}),
    .mi({open_n1765,mem_la_wdata[7]}),
    .f({_al_u1109_o,n17[7]}),
    .q({open_n1781,\uart/uart_odr [7]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("A*~B*C*~D+A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b1110111010100000),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b1110111011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1110|uart/reg3_b2  (
    .a({\uart/uart_status_txd [1],_al_u826_o}),
    .b({\uart/uart_odr [3],_al_u827_o}),
    .c({\uart/uart_odr [4],_al_u828_o}),
    .ce(\uart/mux15_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\uart/uart_status_txd [0],\picorv32_core/pcpi_rs1$2$ }),
    .e({\uart/uart_odr [2],mem_la_wdata[2]}),
    .mi({open_n1783,mem_la_wdata[2]}),
    .f({_al_u1110_o,_al_u851_o}),
    .q({open_n1799,\uart/uart_odr [2]}));  // ../src/uart.v(102)
  // ../src/uart.v(145)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~C*D*~B))"),
    //.LUT1("(~C*~(A*~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100010101010),
    .INIT_LUT1(16'b0000111100000111),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1112|uart/txd_o_reg  (
    .a({txd_pad,_al_u1109_o}),
    .b({_al_u799_o,_al_u1111_o}),
    .c({\uart/uart_status_txd [3],_al_u1113_o}),
    .ce(\uart/n30 ),
    .clk(clk_pad),
    .d({\uart/uart_status_txd [0],_al_u1112_o}),
    .sr(resetn_placeOpt_1),
    .f({_al_u1112_o,open_n1812}),
    .q({open_n1816,txd_pad}));  // ../src/uart.v(145)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("~A*D*C*B"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("~A*~D*~C*B+~A*D*~C*B+~A*D*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b0100000000000000),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b0100010000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1113|uart/reg3_b1  (
    .a({\uart/uart_status_txd [2],_al_u826_o}),
    .b({\uart/uart_status_txd [1],_al_u827_o}),
    .c({\uart/uart_status_txd [0],_al_u828_o}),
    .ce(\uart/mux15_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\uart/uart_odr [1],\picorv32_core/pcpi_rs1$1$ }),
    .e({\uart/uart_odr [0],mem_la_wdata[1]}),
    .mi({open_n1818,mem_la_wdata[1]}),
    .f({_al_u1113_o,_al_u829_o}),
    .q({open_n1834,\uart/uart_odr [1]}));  // ../src/uart.v(102)
  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C))"),
    //.LUT1("(~D*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000010001010),
    .INIT_LUT1(16'b0000000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1116|picorv32_core/reg1_b0  (
    .a({\picorv32_core/mem_xfer_placeOpt_1 ,resetn_placeOpt_13}),
    .b({\picorv32_core/mem_state [0],\picorv32_core/mem_state [0]}),
    .c({open_n1835,trap_pad}),
    .clk(clk_pad),
    .d({\picorv32_core/mem_state [1],_al_u1619_o}),
    .f({\picorv32_core/mux59_sel_is_5_o ,open_n1850}),
    .q({open_n1854,\picorv32_core/mem_state [0]}));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(~C)"),
    //.LUT1("(~B*~D)"),
    .INIT_LUT0(16'b0000111100001111),
    .INIT_LUT1(16'b0000000000110011),
    .MODE("LOGIC"))
    \_al_u1117|_al_u2481  (
    .b({\picorv32_core/n30 [10],open_n1857}),
    .c({open_n1858,\picorv32_core/compressed_instr }),
    .d({\picorv32_core/n30 [11],open_n1861}),
    .f({_al_u1117_o,\picorv32_core/n501 [2]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~A*~B*~D*~C+~A*~B*~D*C"),
    //.LUTG0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0101010001010100),
    .INIT_LUTF1(16'b0000000000010001),
    .INIT_LUTG0(16'b0101000001010000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1118|_al_u2227  (
    .a({\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/pcpi_rs1$12$ }),
    .b({\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .c({open_n1880,\picorv32_core/mem_do_wdata }),
    .d({\picorv32_core/pcpi_rs1$17$ ,open_n1883}),
    .e({\picorv32_core/pcpi_rs1$21$ ,_al_u1546_o_placeOpt_7}),
    .f({_al_u1118_o,_al_u2227_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((~B*~C*D)*~(A)*~(0)+(~B*~C*D)*A*~(0)+~((~B*~C*D))*A*0+(~B*~C*D)*A*0)"),
    //.LUT1("~((~B*~C*D)*~(A)*~(1)+(~B*~C*D)*A*~(1)+~((~B*~C*D))*A*1+(~B*~C*D)*A*1)"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b0101010101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1119 (
    .a({_al_u1118_o,_al_u1118_o}),
    .b({\picorv32_core/n30 [15],\picorv32_core/n30 [15]}),
    .c({\picorv32_core/n30 [19],\picorv32_core/n30 [19]}),
    .d({_al_u1117_o,_al_u1117_o}),
    .mi({open_n1916,_al_u700_o}),
    .fx({open_n1921,_al_u1119_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*~(B*~D)))"),
    //.LUT1("(~C*~B*~D*~A)"),
    .INIT_LUT0(16'b0101000001010100),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u1120|_al_u2183  (
    .a({\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/pcpi_rs1$16$ }),
    .b({\picorv32_core/pcpi_rs1$19$ ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .c({\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/mem_do_wdata }),
    .d({\picorv32_core/pcpi_rs1$18$ ,_al_u1546_o_placeOpt_2}),
    .f({_al_u1120_o,_al_u2183_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*A)"),
    //.LUT1("(~B*~D*C*A)"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"))
    \_al_u1121|_al_u1493  (
    .a({_al_u1120_o,_al_u700_o_placeOpt_1}),
    .b({\picorv32_core/pcpi_rs1$15$ ,open_n1944}),
    .c({_al_u700_o_placeOpt_1,open_n1945}),
    .d({\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/mem_do_rdata }),
    .f({_al_u1121_o,_al_u1493_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D)"),
    //.LUT1("(~B*~D*~A)"),
    .INIT_LUT0(16'b1111000010101010),
    .INIT_LUT1(16'b0000000000010001),
    .MODE("LOGIC"))
    \_al_u1122|_al_u702  (
    .a({\picorv32_core/n30 [13],\picorv32_core/n30 [6]}),
    .b({_al_u700_o,open_n1966}),
    .c({open_n1967,\picorv32_core/pcpi_rs1$8$ }),
    .d({\picorv32_core/n30 [12],_al_u700_o}),
    .f({_al_u1122_o,mem_la_addr[8]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*B*~C*~(~0*~A))"),
    //.LUTF1("A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(D*B*~C*~(~1*~A))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b1110111011101110),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1124|_al_u1179  (
    .a({_al_u1123_o,_al_u1123_o}),
    .b({_al_u1121_o,_al_u1172_o}),
    .c({open_n1988,_al_u1119_o}),
    .d({open_n1991,_al_u1173_o}),
    .e({_al_u1119_o,_al_u1121_o}),
    .f({_al_u1124_o,_al_u1179_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((~C*~D)*~((~0*~A))*~(B)+(~C*~D)*(~0*~A)*~(B)+~((~C*~D))*(~0*~A)*B+(~C*~D)*(~0*~A)*B)"),
    //.LUT1("~((~C*~D)*~((~1*~B))*~(A)+(~C*~D)*(~1*~B)*~(A)+~((~C*~D))*(~1*~B)*A+(~C*~D)*(~1*~B)*A)"),
    .INIT_LUT0(16'b1011101110111000),
    .INIT_LUT1(16'b1111111111111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1125 (
    .a({_al_u700_o_placeOpt_1,\picorv32_core/pcpi_rs1$25$ }),
    .b({\picorv32_core/pcpi_rs1$25$ ,_al_u700_o_placeOpt_1}),
    .c({\picorv32_core/n30 [23],\picorv32_core/n30 [23]}),
    .d({\picorv32_core/n30 [24],\picorv32_core/n30 [24]}),
    .mi({open_n2024,\picorv32_core/pcpi_rs1$26$ }),
    .fx({open_n2029,\eq1/or_xor_i0$13$_i1$13$_o_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("A*~C*B*~D+A*C*B*~D+A*~C*B*D+A*C*B*D"),
    //.LUTG0("~B*A*~C*D+B*A*~C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG1("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1010101000000000),
    .INIT_LUTG1(16'b1101110111011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1126|_al_u1749  (
    .a({_al_u700_o_placeOpt_1,_al_u1313_o}),
    .b({\picorv32_core/pcpi_rs1$28$ ,open_n2032}),
    .d({open_n2037,\picorv32_core/n667_lutinv }),
    .e({\picorv32_core/n30 [26],\picorv32_core/pcpi_rs1$28$ }),
    .f({_al_u1126_o,\picorv32_core/sel43_b28/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0101010001010100),
    .INIT_LUTF1(16'b0101010100110011),
    .INIT_LUTG0(16'b0101000001010000),
    .INIT_LUTG1(16'b0101010100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1127|_al_u2052  (
    .a({\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/pcpi_rs1$27$ }),
    .b({\picorv32_core/n30 [25],\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .c({open_n2058,\picorv32_core/mem_do_wdata }),
    .d({_al_u700_o_placeOpt_1,open_n2061}),
    .e({open_n2062,_al_u1546_o_placeOpt_1}),
    .f({_al_u1127_o,_al_u2052_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("A*~B*C*~D+A*~B*C*D"),
    //.LUTG0("~A*B*~C*~D+A*B*~C*~D"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0010000000100000),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1129|_al_u1168  (
    .a({_al_u1128_o,open_n2083}),
    .b({_al_u1126_o,_al_u1126_o}),
    .c({_al_u1127_o,\eq1/or_xor_i0$13$_i1$13$_o_lutinv }),
    .d({open_n2086,\eq1/or_xor_i0$17$_i1$17$_o_lutinv }),
    .e({\eq1/or_xor_i0$13$_i1$13$_o_lutinv ,_al_u1127_o}),
    .f({_al_u1129_o,_al_u1168_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*~(B*~D)))"),
    //.LUT1("(~A*~D*~C)"),
    .INIT_LUT0(16'b0101000001010100),
    .INIT_LUT1(16'b0000000000000101),
    .MODE("LOGIC"))
    \_al_u1130|_al_u2032  (
    .a({\picorv32_core/pcpi_rs1$31$ ,\picorv32_core/pcpi_rs1$29$ }),
    .b({open_n2107,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .c({\picorv32_core/pcpi_rs1$29$ ,\picorv32_core/mem_do_wdata }),
    .d({\picorv32_core/pcpi_rs1$30$ ,_al_u1546_o_placeOpt_7}),
    .f({_al_u1130_o,_al_u2032_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((~A*~D*~C)*~(B)*~(0)+(~A*~D*~C)*B*~(0)+~((~A*~D*~C))*B*0+(~A*~D*~C)*B*0)"),
    //.LUT1("~((~A*~D*~C)*~(B)*~(1)+(~A*~D*~C)*B*~(1)+~((~A*~D*~C))*B*1+(~A*~D*~C)*B*1)"),
    .INIT_LUT0(16'b1111111111111010),
    .INIT_LUT1(16'b0011001100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1131 (
    .a({\picorv32_core/n30 [27],\picorv32_core/n30 [27]}),
    .b({_al_u1130_o,_al_u1130_o}),
    .c({\picorv32_core/n30 [29],\picorv32_core/n30 [29]}),
    .d({\picorv32_core/n30 [28],\picorv32_core/n30 [28]}),
    .mi({open_n2140,_al_u700_o_placeOpt_1}),
    .fx({open_n2145,\eq1/or_xor_i0$17$_i1$17$_o_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~C*~B*~D)*~(A)*~(0)+(~C*~B*~D)*A*~(0)+~((~C*~B*~D))*A*0+(~C*~B*~D)*A*0)"),
    //.LUTF1("~B*~D*~C*~A+B*~D*~C*~A+~B*~D*C*~A+B*~D*C*~A"),
    //.LUTG0("~((~C*~B*~D)*~(A)*~(1)+(~C*~B*~D)*A*~(1)+~((~C*~B*~D))*A*1+(~C*~B*~D)*A*1)"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1111111111111100),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b0101010101010101),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1132|_al_u1133  (
    .a({\picorv32_core/pcpi_rs1$23$ ,_al_u1132_o}),
    .b({open_n2148,\picorv32_core/n30 [21]}),
    .c({open_n2149,\picorv32_core/n30 [20]}),
    .d({\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/n30 [22]}),
    .e({\picorv32_core/pcpi_rs1$24$ ,_al_u700_o}),
    .f({_al_u1132_o,_al_u1133_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*A*~C*~B+~D*~A*C*~B+~D*A*C*~B+~D*A*~C*B+~D*~A*C*B+~D*A*C*B"),
    //.LUTF1("~A*B*~D*~C+A*B*~D*~C+~A*B*D*~C+A*B*D*~C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG0("~D*~A*C*~B+~D*A*C*~B+~D*~A*C*B+~D*A*C*B"),
    //.LUTG1("A*B*~D*~C+A*B*D*~C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    .INIT_LUTF0(16'b0000000011111010),
    .INIT_LUTF1(16'b1110110011101100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1110100011101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1134|_al_u2140  (
    .a({\picorv32_core/mem_wordsize [0],\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .b({\picorv32_core/mem_wordsize [1],open_n2172}),
    .c({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/mem_do_wdata }),
    .d({open_n2175,\picorv32_core/pcpi_rs1$1$ }),
    .e({\picorv32_core/pcpi_rs1$0$ ,_al_u1546_o_placeOpt_1}),
    .f({_al_u1134_o,_al_u2140_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~A*~B*C*D)"),
    //.LUTF1("(~0*~A*~B*C*D)"),
    //.LUTG0("(~1*~A*~B*C*D)"),
    //.LUTG1("(~1*~A*~B*C*D)"),
    .INIT_LUTF0(16'b0001000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1135|_al_u1137  (
    .a({_al_u1133_o,_al_u1133_o}),
    .b({\eq1/or_xor_i0$17$_i1$17$_o_lutinv ,\eq1/or_xor_i0$17$_i1$17$_o_lutinv }),
    .c({_al_u1129_o,_al_u1129_o}),
    .d({_al_u1124_o,_al_u1124_o}),
    .e({_al_u1134_o,_al_u1136_o}),
    .f({n9,n7}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*~(B*~D)))"),
    //.LUT1("(A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUT0(16'b0101000001010100),
    .INIT_LUT1(16'b1110111011001000),
    .MODE("LOGIC"))
    \_al_u1136|_al_u2260  (
    .a({\picorv32_core/mem_wordsize [0],\picorv32_core/pcpi_rs1$0$ }),
    .b({\picorv32_core/mem_wordsize [1],\picorv32_core/mem_do_prefetch_placeOpt_8 }),
    .c({\picorv32_core/pcpi_rs1$0$ ,\picorv32_core/mem_do_wdata }),
    .d({\picorv32_core/pcpi_rs1$1$ ,_al_u1546_o_placeOpt_8}),
    .f({_al_u1136_o,_al_u2260_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*D+~A*B*~C*D+A*~B*C*D+~A*B*C*D"),
    //.LUTF1("A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("A*~B*~C*D+A*~B*C*D"),
    //.LUTG1("A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*B*~C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0110011000000000),
    .INIT_LUTF1(16'b1100110011101110),
    .INIT_LUTG0(16'b0010001000000000),
    .INIT_LUTG1(16'b1000100011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1138|_al_u1660  (
    .a({\picorv32_core/mem_wordsize [0],\picorv32_core/mem_wordsize [0]}),
    .b({\picorv32_core/mem_wordsize [1],\picorv32_core/mem_wordsize [1]}),
    .d({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$1$ }),
    .e({\picorv32_core/pcpi_rs1$0$ ,\picorv32_core/pcpi_rs1$0$ }),
    .f({_al_u1138_o,_al_u1660_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~A*~B*C*D)"),
    //.LUT1("(~1*~A*~B*D*C)"),
    .INIT_LUT0(16'b0001000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1139 (
    .a({_al_u1133_o,_al_u1133_o}),
    .b({\eq1/or_xor_i0$17$_i1$17$_o_lutinv ,\eq1/or_xor_i0$17$_i1$17$_o_lutinv }),
    .c({_al_u1124_o,_al_u1129_o}),
    .d({_al_u1129_o,_al_u1124_o}),
    .mi({open_n2274,_al_u1138_o}),
    .fx({open_n2279,n13}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~A*~B*C*D)"),
    //.LUT1("(~1*~A*~B*D*C)"),
    .INIT_LUT0(16'b0001000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1141 (
    .a({_al_u1133_o,_al_u1133_o}),
    .b({\eq1/or_xor_i0$17$_i1$17$_o_lutinv ,\eq1/or_xor_i0$17$_i1$17$_o_lutinv }),
    .c({_al_u1124_o,_al_u1129_o}),
    .d({_al_u1129_o,_al_u1124_o}),
    .mi({open_n2294,_al_u1140_o}),
    .fx({open_n2299,n11}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*~C*~B*A)"),
    //.LUTF1("(~0*~D*~C*B*A)"),
    //.LUTG0("(1*~D*~C*~B*A)"),
    //.LUTG1("(~1*~D*~C*B*A)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1143|_al_u1092  (
    .a({\picorv32_core/n328_lutinv ,_al_u1091_o}),
    .b({_al_u1091_o,\picorv32_core/mem_rdata_q [17]}),
    .c({\picorv32_core/mem_rdata_q [17],\picorv32_core/mem_rdata_q [18]}),
    .d({\picorv32_core/mem_rdata_q [18],\picorv32_core/mem_rdata_q [20]}),
    .e({\picorv32_core/mem_rdata_q [21],\picorv32_core/mem_rdata_q [21]}),
    .f({_al_u1143_o,_al_u1092_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*C*~D"),
    //.LUTF1("(~C*A*(B*~(D)*~(0)+~(B)*D*~(0)+~(B)*~(D)*0))"),
    //.LUTG0("0"),
    //.LUTG1("(~C*A*(B*~(D)*~(1)+~(B)*D*~(1)+~(B)*~(D)*1))"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b0000001000001000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1146|_al_u1287  (
    .a({_al_u982_o,_al_u982_o}),
    .b({1'b0,\picorv32_core/cpu_state [7]}),
    .c(\picorv32_core/cpu_state [6:5]),
    .d({\picorv32_core/cpu_state [5],1'b0}),
    .e(\picorv32_core/cpu_state [7:6]),
    .f({\picorv32_core/n746_lutinv ,\picorv32_core/n664_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("A*B*~C*~D"),
    //.LUTF1("A*~B*C*~D+A*~B*~C*D"),
    //.LUTG0("0"),
    //.LUTG1("A*~B*~C*~D"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000001000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1146|_al_u1287_placeOpt_1  (
    .a({_al_u982_o,_al_u982_o}),
    .b(\picorv32_core/cpu_state [6:5]),
    .c({\picorv32_core/cpu_state [7],\picorv32_core/cpu_state [7]}),
    .d({\picorv32_core/cpu_state [5],\picorv32_core/cpu_state [6]}),
    .e(2'b00),
    .f({open_n2363,\picorv32_core/n664_lutinv_placeOpt_1 }));
  EG_PHY_LSLICE #(
    //.LUTF0("A*B*~C*~D"),
    //.LUTF1("A*~B*C*~D+A*~B*~C*D"),
    //.LUTG0("0"),
    //.LUTG1("A*~B*~C*~D"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000001000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1146|_al_u1287_placeOpt_2  (
    .a({_al_u982_o,_al_u982_o}),
    .b(\picorv32_core/cpu_state [6:5]),
    .c({\picorv32_core/cpu_state [7],\picorv32_core/cpu_state [7]}),
    .d({\picorv32_core/cpu_state [5],1'b0}),
    .e({1'b0,\picorv32_core/cpu_state [6]}),
    .f({open_n2386,\picorv32_core/n664_lutinv_placeOpt_2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*C*~D"),
    //.LUTF1("A*B*~C*~D+A*~B*C*~D+A*~B*~C*D"),
    //.LUTG0("0"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b0000001000101000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1146|_al_u1287_placeOpt_3  (
    .a({_al_u982_o,_al_u982_o}),
    .b({1'b0,\picorv32_core/cpu_state [7]}),
    .c({\picorv32_core/cpu_state [5],\picorv32_core/cpu_state [5]}),
    .d({\picorv32_core/cpu_state [7],1'b0}),
    .e({\picorv32_core/cpu_state [6],\picorv32_core/cpu_state [6]}),
    .f({open_n2409,\picorv32_core/n664_lutinv_placeOpt_3 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*C*~D"),
    //.LUTF1("~A*B*C*~D+~A*B*~C*D"),
    //.LUTG0("0"),
    //.LUTG1("~A*B*~C*~D"),
    .INIT_LUTF0(16'b0000000001000000),
    .INIT_LUTF1(16'b0000010001000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1146|_al_u1287_placeOpt_4  (
    .a({\picorv32_core/cpu_state [6],\picorv32_core/cpu_state [7]}),
    .b({_al_u982_o,_al_u982_o}),
    .c({\picorv32_core/cpu_state [5],\picorv32_core/cpu_state [5]}),
    .d({\picorv32_core/cpu_state [7],1'b0}),
    .e({1'b0,\picorv32_core/cpu_state [6]}),
    .f({open_n2432,\picorv32_core/n664_lutinv_placeOpt_4 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*C*~D"),
    //.LUTF1("~A*B*C*~D+~A*B*~C*D"),
    //.LUTG0("0"),
    //.LUTG1("~A*B*~C*~D"),
    .INIT_LUTF0(16'b0000000001000000),
    .INIT_LUTF1(16'b0000010001000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1146|_al_u1287_placeOpt_5  (
    .a({\picorv32_core/cpu_state [6],\picorv32_core/cpu_state [7]}),
    .b({_al_u982_o,_al_u982_o}),
    .c({\picorv32_core/cpu_state [5],\picorv32_core/cpu_state [5]}),
    .d(\picorv32_core/cpu_state [7:6]),
    .e(2'b00),
    .f({open_n2455,\picorv32_core/n664_lutinv_placeOpt_5 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~A*C*~B*D)"),
    //.LUTF1("A*~B*~C*D+~A*~B*C*D"),
    //.LUTG0("(~1*~A*C*~B*D)"),
    //.LUTG1("~A*~B*~C*D"),
    .INIT_LUTF0(16'b0001000000000000),
    .INIT_LUTF1(16'b0001001000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1146|_al_u1287_placeOpt_6  (
    .a(\picorv32_core/cpu_state [7:6]),
    .b({\picorv32_core/cpu_state [6],1'b0}),
    .c({\picorv32_core/cpu_state [5],\picorv32_core/cpu_state [5]}),
    .d({_al_u982_o,_al_u982_o}),
    .e({1'b0,\picorv32_core/cpu_state [7]}),
    .f({open_n2478,\picorv32_core/n664_lutinv_placeOpt_6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*C*~A*B)"),
    //.LUTF1("(~B*D*(A*~(C)*~(0)+~(A)*C*~(0)+~(A)*~(C)*0))"),
    //.LUTG0("(~1*~D*C*~A*B)"),
    //.LUTG1("(~B*D*(A*~(C)*~(1)+~(A)*C*~(1)+~(A)*~(C)*1))"),
    .INIT_LUTF0(16'b0000000001000000),
    .INIT_LUTF1(16'b0001001000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1146|_al_u1287_placeOpt_7  (
    .a(2'b00),
    .b({\picorv32_core/cpu_state [6],_al_u982_o}),
    .c({\picorv32_core/cpu_state [5],\picorv32_core/cpu_state [5]}),
    .d({_al_u982_o,\picorv32_core/cpu_state [6]}),
    .e({\picorv32_core/cpu_state [7],\picorv32_core/cpu_state [7]}),
    .f({open_n2501,\picorv32_core/n664_lutinv_placeOpt_7 }));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG0("~D*B*~C*A+D*B*~C*A"),
    //.LUTG1("~A*~B*~C*D+~A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000100000000),
    .INIT_LUTG0(16'b0000100000001000),
    .INIT_LUTG1(16'b0001000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1147|picorv32_core/trap_reg  (
    .a({\picorv32_core/cpu_state [6],\picorv32_core/cpu_state [7]}),
    .b({\picorv32_core/cpu_state [7],_al_u980_o}),
    .c({open_n2507,\picorv32_core/cpu_state [6]}),
    .clk(clk_pad),
    .d({_al_u980_o,open_n2509}),
    .e({open_n2510,_al_u982_o}),
    .sr(resetn_placeOpt_8),
    .f({_al_u1147_o,\picorv32_core/n662 }),
    .q({open_n2528,trap_pad}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*~C*~B*A)"),
    //.LUTF1("(~0*~B*A*~D*C)"),
    //.LUTG0("(~1*D*~C*~B*A)"),
    //.LUTG1("(~1*~B*A*~D*C)"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b0000000000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1148|_al_u1150  (
    .a({\picorv32_core/cpu_state [1],_al_u1147_o}),
    .b({\picorv32_core/cpu_state [2],\picorv32_core/cpu_state [0]}),
    .c({_al_u1147_o,\picorv32_core/cpu_state [1]}),
    .d({\picorv32_core/cpu_state [0],\picorv32_core/cpu_state [2]}),
    .e({\picorv32_core/cpu_state [3],\picorv32_core/cpu_state [3]}),
    .f({\picorv32_core/n668_lutinv ,\picorv32_core/n667_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*B*A)"),
    //.LUT1("(~1*~C*~D*A*B)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1149 (
    .a({\picorv32_core/cpu_state [0],_al_u1147_o}),
    .b({_al_u1147_o,\picorv32_core/cpu_state [0]}),
    .c(\picorv32_core/cpu_state [2:1]),
    .d({\picorv32_core/cpu_state [1],\picorv32_core/cpu_state [2]}),
    .mi({open_n2563,\picorv32_core/cpu_state [3]}),
    .fx({open_n2568,\picorv32_core/n669_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*B*A)"),
    //.LUT1("(~1*~D*~C*B*A)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1149_placeOpt_1 (
    .a({_al_u1147_o,_al_u1147_o}),
    .b({\picorv32_core/cpu_state [0],\picorv32_core/cpu_state [0]}),
    .c({\picorv32_core/cpu_state [1],\picorv32_core/cpu_state [1]}),
    .d({\picorv32_core/cpu_state [2],\picorv32_core/cpu_state [2]}),
    .mi({open_n2583,\picorv32_core/cpu_state [3]}),
    .fx({open_n2588,\picorv32_core/n669_lutinv_placeOpt_1 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*B*A)"),
    //.LUT1("(~1*~D*~C*B*A)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1149_placeOpt_2 (
    .a({_al_u1147_o,_al_u1147_o}),
    .b({\picorv32_core/cpu_state [0],\picorv32_core/cpu_state [0]}),
    .c({\picorv32_core/cpu_state [1],\picorv32_core/cpu_state [1]}),
    .d({\picorv32_core/cpu_state [2],\picorv32_core/cpu_state [2]}),
    .mi({open_n2603,\picorv32_core/cpu_state [3]}),
    .fx({open_n2608,\picorv32_core/n669_lutinv_placeOpt_2 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*B*A)"),
    //.LUT1("(~1*~C*~D*A*B)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1149_placeOpt_3 (
    .a({\picorv32_core/cpu_state [0],_al_u1147_o}),
    .b({_al_u1147_o,\picorv32_core/cpu_state [0]}),
    .c(\picorv32_core/cpu_state [2:1]),
    .d({\picorv32_core/cpu_state [1],\picorv32_core/cpu_state [2]}),
    .mi({open_n2623,\picorv32_core/cpu_state [3]}),
    .fx({open_n2628,\picorv32_core/n669_lutinv_placeOpt_3 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*B*A)"),
    //.LUT1("(~1*~D*~C*B*A)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1149_placeOpt_4 (
    .a({_al_u1147_o,_al_u1147_o}),
    .b({\picorv32_core/cpu_state [0],\picorv32_core/cpu_state [0]}),
    .c({\picorv32_core/cpu_state [1],\picorv32_core/cpu_state [1]}),
    .d({\picorv32_core/cpu_state [2],\picorv32_core/cpu_state [2]}),
    .mi({open_n2643,\picorv32_core/cpu_state [3]}),
    .fx({open_n2648,\picorv32_core/n669_lutinv_placeOpt_4 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*B*~(C*~(0*~D)))"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D"),
    //.LUTG0("(~A*B*~(C*~(1*~D)))"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000010000000100),
    .INIT_LUTF1(16'b0000000010101010),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1153|_al_u1906  (
    .a({_al_u1151_o,\picorv32_core/n663 }),
    .b({open_n2651,_al_u1151_o}),
    .c({open_n2652,\picorv32_core/n666_lutinv }),
    .d({\picorv32_core/n666_lutinv ,_al_u1216_o}),
    .e({\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ,\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .f({_al_u1153_o,_al_u1906_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*(A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D))"),
    //.LUTF1("0"),
    //.LUTG0("(~1*(A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D))"),
    //.LUTG1("~A*~B*~C*D+~A*B*~C*D"),
    .INIT_LUTF0(16'b0000011111111110),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1159|_al_u1072  (
    .a({\uart/uart_status_rxd [0],\uart/uart_status_rxd [0]}),
    .b({open_n2675,\uart/uart_status_rxd [1]}),
    .c({\uart/uart_status_rxd [2],\uart/uart_status_rxd [2]}),
    .d({\uart/uart_status_rxd [3],\uart/uart_status_rxd [3]}),
    .e({\uart/uart_status_rxd [1],\uart/uart_cnt_rx [0]}),
    .f({_al_u1159_o,_al_u1072_o}));
  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*~B*A)"),
    //.LUT1("(D*~(~A*B*~C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000100000),
    .INIT_LUT1(16'b1111101100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1160|uart/uart_status_rx_reg  (
    .a({\uart/uart_cnt_rx [2],_al_u1063_o}),
    .b(\uart/uart_cnt_rx [1:0]),
    .c({\uart/uart_cnt_rx [0],\uart/uart_cnt_rx [1]}),
    .ce(\picorv32_core/n524$4$_en ),
    .clk(clk_pad),
    .d({_al_u1159_o,\uart/uart_cnt_rx [2]}),
    .sr(resetn_placeOpt_9),
    .f({_al_u1160_o,\uart/mux51_b0_sel_is_3_o }),
    .q({open_n2713,\uart/uart_status_rx }));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(C)*~(D)*~((~0*B))+A*~(C)*~(D)*~((~0*B))+~(A)*C*~(D)*~((~0*B))+~(A)*C*D*~((~0*B))+~(A)*C*D*(~0*B))"),
    //.LUT1("(~(A)*~(C)*~(D)*~((~1*B))+A*~(C)*~(D)*~((~1*B))+~(A)*C*~(D)*~((~1*B))+~(A)*C*D*~((~1*B))+~(A)*C*D*(~1*B))"),
    .INIT_LUT0(16'b0101000000010011),
    .INIT_LUT1(16'b0101000001011111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1164 (
    .a({\uart/n77 [0],\uart/n77 [0]}),
    .b({_al_u1070_o,_al_u1070_o}),
    .c({\uart/n51_lutinv ,\uart/n51_lutinv }),
    .d({\uart/uart_status_rxd [0],\uart/uart_status_rxd [0]}),
    .mi({open_n2726,rxd_pad}),
    .fx({open_n2731,_al_u1164_o}));
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(~B*~(A*D*C)))"),
    //.LUTF1("(~A*B)"),
    //.LUTG0("(1*~(~B*~(A*D*C)))"),
    //.LUTG1("(~A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0100010001000100),
    .INIT_LUTG0(16'b1110110011001100),
    .INIT_LUTG1(16'b0100010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1167|picorv32_core/mem_la_secondword_reg  (
    .a({\picorv32_core/n111 ,\picorv32_core/mem_la_firstword_xfer }),
    .b({\picorv32_core/mux59_sel_is_5_o ,\picorv32_core/n25 }),
    .c({open_n2734,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .ce(\picorv32_core/mux59_sel_is_5_o ),
    .clk(clk_pad),
    .d({open_n2735,\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }),
    .e({open_n2736,resetn_placeOpt_15}),
    .sr(\picorv32_core/n111 ),
    .f({\picorv32_core/mux68_b0_sel_is_2_o ,\picorv32_core/mem_la_read }),
    .q({open_n2754,\picorv32_core/mem_la_secondword }));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("~((~C*~D)*~((~0*~A))*~(B)+(~C*~D)*(~0*~A)*~(B)+~((~C*~D))*(~0*~A)*B+(~C*~D)*(~0*~A)*B)"),
    //.LUT1("~((~C*~D)*~((~1*~A))*~(B)+(~C*~D)*(~1*~A)*~(B)+~((~C*~D))*(~1*~A)*B+(~C*~D)*(~1*~A)*B)"),
    .INIT_LUT0(16'b1011101110111000),
    .INIT_LUT1(16'b1111111111111100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1169 (
    .a({\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$10$ }),
    .b({_al_u700_o,_al_u700_o}),
    .c({\picorv32_core/n30 [7],\picorv32_core/n30 [7]}),
    .d({\picorv32_core/n30 [8],\picorv32_core/n30 [8]}),
    .mi({open_n2767,\picorv32_core/pcpi_rs1$9$ }),
    .fx({open_n2772,\eq2/or_xor_i0$5$_i1$5$_o_o_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*A*B*D*C)"),
    //.LUTF1("~D*~B*~A*~C+~D*~B*A*~C"),
    //.LUTG0("(1*A*B*D*C)"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1170|_al_u1174  (
    .a({open_n2775,_al_u1172_o}),
    .b({\eq2/or_xor_i0$5$_i1$5$_o_o_lutinv ,_al_u1170_o}),
    .c({mem_la_addr[4],_al_u1124_o}),
    .d({mem_la_addr[11],_al_u1168_o}),
    .e({_al_u1133_o,_al_u1173_o}),
    .f({_al_u1170_o,n16}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D*~(B*~(0)*~(A)+B*0*~(A)+~(B)*0*A+B*0*A))"),
    //.LUT1("(~C*~D*~(B*~(1)*~(A)+B*1*~(A)+~(B)*1*A+B*1*A))"),
    .INIT_LUT0(16'b0000000000001011),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1172 (
    .a({_al_u700_o,_al_u700_o}),
    .b({\picorv32_core/n30 [6],\picorv32_core/n30 [6]}),
    .c({mem_la_addr[7],mem_la_addr[7]}),
    .d({\eq2/or_xor_i0$1$_i1$1$_o_o_lutinv ,\eq2/or_xor_i0$1$_i1$1$_o_o_lutinv }),
    .mi({open_n2810,\picorv32_core/pcpi_rs1$8$ }),
    .fx({open_n2815,_al_u1172_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(B*~A*~D*~C)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("LOGIC"))
    \_al_u1175|_al_u709  (
    .a({mem_la_addr[11],open_n2818}),
    .b({mem_la_addr[4],\picorv32_core/pcpi_rs1$11$ }),
    .c({_al_u1133_o,_al_u700_o}),
    .d({\eq2/or_xor_i0$5$_i1$5$_o_o_lutinv ,\picorv32_core/n30 [9]}),
    .f({_al_u1175_o,mem_la_addr[11]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~D)"),
    //.LUT1("(A*D*C)"),
    .INIT_LUT0(16'b0000000001010000),
    .INIT_LUT1(16'b1010000000000000),
    .MODE("LOGIC"))
    \_al_u1176|_al_u1173  (
    .a({_al_u1128_o,mem_la_addr[2]}),
    .c({mem_la_addr[3],_al_u1128_o}),
    .d({mem_la_addr[2],mem_la_addr[3]}),
    .f({\uart/u7_sel_is_3_o ,_al_u1173_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*C*B*A*D)"),
    //.LUT1("(~1*C*B*A*D)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1178 (
    .a({_al_u1168_o,_al_u1168_o}),
    .b({_al_u1175_o,_al_u1175_o}),
    .c({_al_u1172_o,_al_u1172_o}),
    .d({_al_u1124_o,_al_u1124_o}),
    .mi({open_n2873,_al_u1128_o}),
    .fx({open_n2878,\uart/mux14_b0_sel_is_1_o }));
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(B*~C)"),
    //.LUTG0("C*D*A*B"),
    //.LUTG1("(B*~C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000110000001100),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1181|uart/reg2_b0  (
    .a({open_n2881,_al_u1175_o}),
    .b({_al_u1128_o,_al_u1172_o}),
    .c({_al_u812_o,\uart/mux9_b0_sel_is_3_o }),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({open_n2882,_al_u1168_o}),
    .e({open_n2883,_al_u1124_o}),
    .mi({open_n2885,mem_la_wdata[0]}),
    .sr(resetn),
    .f({\uart/mux9_b0_sel_is_3_o ,\uart/mux12_b0_sel_is_3_o }),
    .q({open_n2900,\uart/uart_bsrr [0]}));  // ../src/uart.v(102)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~0*~(~D*C))*~(B*A))"),
    //.LUTF1("~B*~A*~D*~C+B*~A*~D*~C+~B*~A*~D*C+B*~A*~D*C"),
    //.LUTG0("(~(~1*~(~D*C))*~(B*A))"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000001110000),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b0111011101110111),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1183|picorv32_core/latched_stalu_reg  (
    .a({\picorv32_core/n666_lutinv ,_al_u1183_o}),
    .b({open_n2901,_al_u1184_o}),
    .c({open_n2902,\picorv32_core/n666_lutinv }),
    .clk(clk_pad),
    .d({\picorv32_core/n667_lutinv ,\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .e({\picorv32_core/n746_lutinv ,\picorv32_core/latched_stalu }),
    .sr(resetn_placeOpt_8),
    .f({_al_u1183_o,open_n2918}),
    .q({open_n2922,\picorv32_core/latched_stalu }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*~A)"),
    //.LUT1("(~C*~A)"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"))
    \_al_u1184|_al_u1151  (
    .a({\picorv32_core/n668_lutinv ,\picorv32_core/n746_lutinv }),
    .b({open_n2923,\picorv32_core/n668_lutinv }),
    .c({\picorv32_core/n669_lutinv_placeOpt_1 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .d({open_n2926,\picorv32_core/n667_lutinv }),
    .f({_al_u1184_o,_al_u1151_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~D*~C+~A*~B*~D*C"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    //.LUTG0("~A*~B*~D*~C+~A*~B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000010001),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0001000100010001),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1186|_al_u2083  (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_rdata }),
    .b({open_n2945,\picorv32_core/n576 [24]}),
    .d({open_n2950,\picorv32_core/mem_do_prefetch_placeOpt_4 }),
    .e({\picorv32_core/mem_do_wdata ,_al_u1546_o_placeOpt_5}),
    .f({_al_u1186_o,_al_u2083_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~A*~(~D*~(0*~B)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("(~C*~A*~(~D*~(1*~B)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0000010100000000),
    .INIT_LUTF1(16'b0101010111111111),
    .INIT_LUTG0(16'b0000010100000001),
    .INIT_LUTG1(16'b0101010101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1188|_al_u1187  (
    .a({resetn_placeOpt_17,_al_u1186_o}),
    .b({open_n2971,\picorv32_core/mem_wordsize [0]}),
    .c({\picorv32_core/mem_do_rinst ,\picorv32_core/mem_wordsize [1]}),
    .d({_al_u1187_o,\picorv32_core/pcpi_rs1$0$ }),
    .e({\picorv32_core/reg_pc [0],\picorv32_core/pcpi_rs1$1$ }),
    .f({\picorv32_core/mux164_b0_sel_is_0_o ,_al_u1187_o}));
  // ../src/uart.v(263)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+A*B*C*D*~(0)+A*B*~(C)*~(D)*0)"),
    //.LUTF1("(~(C)*~(B)*~(A)*~(D)*~(0)+C*~(B)*~(A)*~(D)*~(0)+~(C)*B*~(A)*~(D)*~(0)+C*B*~(A)*~(D)*~(0)+~(C)*B*A*~(D)*~(0)+~(C)*~(B)*~(A)*D*~(0)+C*~(B)*~(A)*D*~(0)+~(C)*B*~(A)*D*~(0)+~(C)*B*A*D*~(0)+~(C)*~(B)*~(A)*~(D)*0+C*~(B)*~(A)*~(D)*0+~(C)*B*~(A)*~(D)*0+~(C)*~(B)*A*~(D)*0+C*~(B)*A*~(D)*0+~(C)*B*A*~(D)*0+C*B*A*~(D)*0+~(C)*~(B)*~(A)*D*0+C*~(B)*~(A)*D*0+~(C)*B*~(A)*D*0+C*B*~(A)*D*0+~(C)*~(B)*A*D*0+C*~(B)*A*D*0+~(C)*B*A*D*0+C*B*A*D*0)"),
    //.LUTG0("(A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+A*B*C*D*~(1)+A*B*~(C)*~(D)*1)"),
    //.LUTG1("(~(C)*~(B)*~(A)*~(D)*~(1)+C*~(B)*~(A)*~(D)*~(1)+~(C)*B*~(A)*~(D)*~(1)+C*B*~(A)*~(D)*~(1)+~(C)*B*A*~(D)*~(1)+~(C)*~(B)*~(A)*D*~(1)+C*~(B)*~(A)*D*~(1)+~(C)*B*~(A)*D*~(1)+~(C)*B*A*D*~(1)+~(C)*~(B)*~(A)*~(D)*1+C*~(B)*~(A)*~(D)*1+~(C)*B*~(A)*~(D)*1+~(C)*~(B)*A*~(D)*1+C*~(B)*A*~(D)*1+~(C)*B*A*~(D)*1+C*B*A*~(D)*1+~(C)*~(B)*~(A)*D*1+C*~(B)*~(A)*D*1+~(C)*B*~(A)*D*1+C*B*~(A)*D*1+~(C)*~(B)*A*D*1+C*~(B)*A*D*1+~(C)*B*A*D*1+C*B*A*D*1)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101110000000),
    .INIT_LUTF1(16'b0001110101011101),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b1111111110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1189|uart/reg5_b2  (
    .a({\uart/uart_status_rxd [1],\uart/n77 [2]}),
    .b({\uart/n51_lutinv ,\uart/n51_lutinv }),
    .c({\uart/n77 [1],\uart/uart_status_rxd [1]}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({\uart/uart_status_rxd [2],\uart/uart_status_rxd [2]}),
    .e({\uart/uart_status_rxd [3],\uart/uart_status_rxd [3]}),
    .sr(resetn_placeOpt_9),
    .f({_al_u1189_o,open_n3008}),
    .q({open_n3012,\uart/uart_status_rxd [2]}));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~A)"),
    //.LUT1("(D*~B)"),
    .INIT_LUT0(16'b0000010100000000),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"))
    \_al_u1190|_al_u1161  (
    .a({open_n3013,\uart/uart_cnt_rx [0]}),
    .b({_al_u1086_o,open_n3014}),
    .c({open_n3015,\uart/uart_cnt_rx [1]}),
    .d({\uart/n51_lutinv ,\uart/uart_cnt_rx [2]}),
    .f({\uart/mux37_b0_sel_is_3_o ,\uart/n51_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~(B*C*A*D))"),
    //.LUT1("~(~1*~(B*C*A*D))"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1192 (
    .a({_al_u1168_o,_al_u1168_o}),
    .b({\uart/n9_lutinv ,\uart/n9_lutinv }),
    .c({_al_u1175_o,_al_u1175_o}),
    .d({_al_u1179_o,_al_u1179_o}),
    .mi({open_n3048,_al_u1076_o}),
    .fx({open_n3053,\picorv32_core/n524$4$_en_al_n602 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("~A*~B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*B*~C*D"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("~A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b0000100100001001),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b1001000010010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1194|_al_u841  (
    .a({\picorv32_core/pcpi_rs2$15$ ,_al_u826_o}),
    .b({\picorv32_core/pcpi_rs1$15$ ,_al_u827_o}),
    .c({\picorv32_core/pcpi_rs2$16$ ,_al_u828_o}),
    .d({open_n3058,\picorv32_core/pcpi_rs1$15$ }),
    .e({\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/pcpi_rs2$15$ }),
    .f({_al_u1194_o,_al_u841_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("D*~B*~C*~A+D*B*~C*A"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("D*~B*C*~A+D*B*C*A"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b0000100100000000),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b1001000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1195|_al_u839  (
    .a({\picorv32_core/pcpi_rs1$14$ ,_al_u826_o}),
    .b({\picorv32_core/pcpi_rs2$14$ ,_al_u827_o}),
    .c({\picorv32_core/pcpi_rs2$13$ ,_al_u828_o}),
    .d({_al_u1194_o,\picorv32_core/pcpi_rs1$14$ }),
    .e({\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/pcpi_rs2$14$ }),
    .f({_al_u1195_o,_al_u839_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*B*~A*~C+~D*~B*A*~C+~D*B*A*~C+~D*B*~A*C+~D*~B*A*C+~D*B*A*C"),
    //.LUTF1("~D*~B*~A*~C+D*B*~A*~C+~D*~B*A*~C+D*B*A*~C"),
    //.LUTG0("~D*~B*A*~C+~D*B*A*~C+~D*~B*A*C+~D*B*A*C"),
    //.LUTG1("~D*~B*~A*C+D*B*~A*C+~D*~B*A*C+D*B*A*C"),
    .INIT_LUTF0(16'b0000000011101110),
    .INIT_LUTF1(16'b0000110000000011),
    .INIT_LUTG0(16'b0000000010101010),
    .INIT_LUTG1(16'b1100000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1196|_al_u2238  (
    .a({open_n3101,\picorv32_core/mem_do_wdata }),
    .b({\picorv32_core/pcpi_rs1$11$ ,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .c({\picorv32_core/pcpi_rs2$12$ ,open_n3102}),
    .d({\picorv32_core/pcpi_rs2$11$ ,\picorv32_core/pcpi_rs1$11$ }),
    .e({\picorv32_core/pcpi_rs1$12$ ,_al_u1546_o_placeOpt_1}),
    .f({_al_u1196_o,_al_u2238_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("D*~B*~C*~A+D*~B*C*A"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("D*B*~C*~A+D*B*C*A"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b0010000100000000),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b1000010000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1197|_al_u831  (
    .a({\picorv32_core/pcpi_rs2$10$ ,_al_u826_o}),
    .b({mem_la_wdata[1],_al_u827_o}),
    .c({\picorv32_core/pcpi_rs1$10$ ,_al_u828_o}),
    .d({_al_u1196_o,\picorv32_core/pcpi_rs1$10$ }),
    .e({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs2$10$ }),
    .f({_al_u1197_o,_al_u831_o}));
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    //.LUT1("(~(A@D)*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100101011001010),
    .INIT_LUT1(16'b1000001001000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1198|uart/reg2_b23  (
    .a({\picorv32_core/pcpi_rs2$23$ ,mem_la_wdata[7]}),
    .b({\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs2$23$ }),
    .c({\picorv32_core/pcpi_rs2$22$ ,\picorv32_core/n734_lutinv }),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\picorv32_core/pcpi_rs1$23$ ,open_n3147}),
    .sr(resetn_placeOpt_12),
    .f({_al_u1198_o,mem_la_wdata[23]}),
    .q({open_n3163,\uart/uart_bsrr [23]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTF1("C*~B*~A*~D+C*B*A*~D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("C*~B*~A*D+C*B*A*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000010010000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1001000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1199|uart/reg2_b21  (
    .a({\picorv32_core/pcpi_rs1$21$ ,open_n3164}),
    .b({\picorv32_core/pcpi_rs2$21$ ,open_n3165}),
    .c({_al_u1198_o,mem_la_wdata[5]}),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\picorv32_core/pcpi_rs2$20$ ,\picorv32_core/n734_lutinv }),
    .e({\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/pcpi_rs2$21$ }),
    .sr(resetn_placeOpt_12),
    .f({_al_u1199_o,mem_la_wdata[21]}),
    .q({open_n3183,\uart/uart_bsrr [21]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    //.LUT1("(~(D@C)*~(B@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101100011011000),
    .INIT_LUT1(16'b1001000000001001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1200|uart/reg2_b19  (
    .a({\picorv32_core/pcpi_rs1$19$ ,\picorv32_core/n734_lutinv }),
    .b({\picorv32_core/pcpi_rs2$19$ ,\picorv32_core/pcpi_rs2$19$ }),
    .c({\picorv32_core/pcpi_rs1$2$ ,mem_la_wdata[3]}),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({mem_la_wdata[2],open_n3184}),
    .sr(resetn_placeOpt_12),
    .f({_al_u1200_o,mem_la_wdata[19]}),
    .q({open_n3200,\uart/uart_bsrr [19]}));  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(0@A)*~(B@D))"),
    //.LUT1("(C*~(1@A)*~(B@D))"),
    .INIT_LUT0(16'b0100000000010000),
    .INIT_LUT1(16'b1000000000100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1201 (
    .a({\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$18$ }),
    .b({\picorv32_core/pcpi_rs2$17$ ,\picorv32_core/pcpi_rs2$17$ }),
    .c({_al_u1200_o,_al_u1200_o}),
    .d({\picorv32_core/pcpi_rs1$17$ ,\picorv32_core/pcpi_rs1$17$ }),
    .mi({open_n3213,\picorv32_core/pcpi_rs2$18$ }),
    .fx({open_n3218,_al_u1201_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*A*D)"),
    //.LUT1("(A*B*C*D)"),
    .INIT_LUT0(16'b1010000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u1202|_al_u1827  (
    .a({_al_u1201_o,\picorv32_core/n734_lutinv }),
    .b({_al_u1199_o,open_n3221}),
    .c({_al_u1197_o,\picorv32_core/latched_is_lu }),
    .d({_al_u1195_o,mem_rdata[18]}),
    .f({_al_u1202_o,\picorv32_core/sel27_b18/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*C*~D+~A*B*~C*D+A*B*C*D"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*C*~D+~A*B*~C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1203|_al_u889  (
    .a({\picorv32_core/pcpi_rs1$9$ ,_al_u826_o}),
    .b({\picorv32_core/pcpi_rs1$0$ ,_al_u827_o}),
    .c({\picorv32_core/pcpi_rs2$9$ ,_al_u828_o}),
    .d({mem_la_wdata[0],\picorv32_core/pcpi_rs1$9$ }),
    .e({open_n3244,\picorv32_core/pcpi_rs2$9$ }),
    .f({_al_u1203_o,_al_u889_o}));
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("D*~B*~C*~A+D*~B*C*A"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("D*B*~C*~A+D*B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b0010000100000000),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b1000010000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1204|uart/reg2_b7  (
    .a({\picorv32_core/pcpi_rs2$8$ ,_al_u826_o}),
    .b({mem_la_wdata[7],_al_u827_o}),
    .c({\picorv32_core/pcpi_rs1$8$ ,_al_u828_o}),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({_al_u1203_o,\picorv32_core/pcpi_rs1$7$ }),
    .e({\picorv32_core/pcpi_rs1$7$ ,mem_la_wdata[7]}),
    .mi({open_n3266,mem_la_wdata[7]}),
    .sr(resetn),
    .f({_al_u1204_o,_al_u885_o}),
    .q({open_n3281,\uart/uart_bsrr [7]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("~A*~D*~C*~B+~A*D*~C*~B+A*~D*C*~B+A*D*C*~B"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("~A*~D*~C*B+~A*D*~C*B+A*~D*C*B+A*D*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b0010000100100001),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b1000010010000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1205|uart/reg2_b6  (
    .a({mem_la_wdata[6],_al_u826_o}),
    .b({mem_la_wdata[5],_al_u827_o}),
    .c({\picorv32_core/pcpi_rs1$6$ ,_al_u828_o}),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({open_n3282,\picorv32_core/pcpi_rs1$6$ }),
    .e({\picorv32_core/pcpi_rs1$5$ ,mem_la_wdata[6]}),
    .mi({open_n3284,mem_la_wdata[6]}),
    .sr(resetn_placeOpt_2),
    .f({_al_u1205_o,_al_u883_o}),
    .q({open_n3299,\uart/uart_bsrr [6]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("0"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("~D*~A*~B*~C+D*~A*B*~C+~D*A*~B*C+D*A*B*C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1206|uart/reg2_b4  (
    .a({\picorv32_core/pcpi_rs1$31$ ,_al_u826_o}),
    .b({\picorv32_core/pcpi_rs1$4$ ,_al_u827_o}),
    .c({\picorv32_core/pcpi_rs2$31$ ,_al_u828_o}),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({mem_la_wdata[4],\picorv32_core/pcpi_rs1$4$ }),
    .e({_al_u1205_o,mem_la_wdata[4]}),
    .mi({open_n3301,mem_la_wdata[4]}),
    .sr(resetn),
    .f({_al_u1206_o,_al_u879_o}),
    .q({open_n3316,\uart/uart_bsrr [4]}));  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTF1("(~(D@B)*~(A@C))"),
    //.LUTG0("0"),
    //.LUTG1("(~(D@B)*~(A@C))"),
    .INIT_LUTF0(16'b1111000011111010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1208|_al_u2011  (
    .a({mem_la_wdata[3],\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .b({\picorv32_core/pcpi_rs1$30$ ,open_n3317}),
    .c({\picorv32_core/pcpi_rs1$3$ ,\picorv32_core/mem_do_wdata }),
    .d({\picorv32_core/pcpi_rs2$30$ ,_al_u1546_o_placeOpt_7}),
    .e({open_n3320,\picorv32_core/pcpi_rs1$30$ }),
    .f({_al_u1208_o,_al_u2011_o}));
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B)*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("A*~B*~C*~D+A*B*C*~D"),
    //.LUTG0("(A*~(B)*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("A*~B*~C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000100100000),
    .INIT_LUTF1(16'b0000000010000010),
    .INIT_LUTG0(16'b0111010101100100),
    .INIT_LUTG1(16'b1000001000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1209|uart/reg2_b29  (
    .a({_al_u1208_o,\picorv32_core/mem_wordsize [0]}),
    .b({\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/mem_wordsize [1]}),
    .c({\picorv32_core/pcpi_rs2$28$ ,\picorv32_core/pcpi_rs2$13$ }),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\picorv32_core/pcpi_rs2$29$ ,\picorv32_core/pcpi_rs2$29$ }),
    .e({\picorv32_core/pcpi_rs1$29$ ,mem_la_wdata[5]}),
    .sr(resetn_placeOpt_12),
    .f({_al_u1209_o,mem_la_wdata[29]}),
    .q({open_n3358,\uart/uart_bsrr [29]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B)*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~A*~B*~D*~C+~A*~B*D*~C+~A*B*~D*C+~A*B*D*C"),
    //.LUTG0("(A*~(B)*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("A*~B*~D*~C+A*~B*D*~C+A*B*~D*C+A*B*D*C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000100100000),
    .INIT_LUTF1(16'b0100000101000001),
    .INIT_LUTG0(16'b0111010101100100),
    .INIT_LUTG1(16'b1000001010000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1210|uart/reg2_b27  (
    .a({\picorv32_core/pcpi_rs2$26$ ,\picorv32_core/mem_wordsize [0]}),
    .b({\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/mem_wordsize [1]}),
    .c({\picorv32_core/pcpi_rs2$27$ ,\picorv32_core/pcpi_rs2$11$ }),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({open_n3359,\picorv32_core/pcpi_rs2$27$ }),
    .e({\picorv32_core/pcpi_rs1$26$ ,mem_la_wdata[3]}),
    .sr(resetn_placeOpt_12),
    .f({_al_u1210_o,mem_la_wdata[27]}),
    .q({open_n3377,\uart/uart_bsrr [27]}));  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(0@C)*~(A@B))"),
    //.LUTF1("0"),
    //.LUTG0("(D*~(1@C)*~(A@B))"),
    //.LUTG1("A*~B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000100100000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1001000000000000),
    .INIT_LUTG1(16'b1010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1212|_al_u1211  (
    .a({_al_u1209_o,\picorv32_core/pcpi_rs2$24$ }),
    .b({open_n3378,\picorv32_core/pcpi_rs1$24$ }),
    .c({_al_u1207_o,\picorv32_core/pcpi_rs1$25$ }),
    .d({_al_u1211_o,_al_u1210_o}),
    .e({_al_u1202_o,\picorv32_core/pcpi_rs2$25$ }),
    .f({\picorv32_core/alu_eq_lutinv ,_al_u1211_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~C*~D*~A*~B+C*~D*~A*~B+~C*~D*A*~B+C*~D*A*~B+~C*~D*~A*B+C*~D*~A*B+~C*~D*A*B+C*~D*A*B"),
    //.LUTG0("B*D*A*~C+B*D*A*C"),
    //.LUTG1("~C*~D*~A*~B+C*~D*~A*~B+~C*D*~A*~B+C*D*~A*~B+~C*~D*~A*B+C*~D*~A*B+~C*D*~A*B+C*D*~A*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b1000100000000000),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1213|picorv32_core/instr_bgeu_reg  (
    .a({\picorv32_core/is_sltiu_bltu_sltu ,\picorv32_core/mem_rdata_q [13]}),
    .b({open_n3401,\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_bgeu ,\picorv32_core/mem_rdata_q [12]}),
    .e({\picorv32_core/alu_ltu ,\picorv32_core/mem_rdata_q [14]}),
    .sr(resetn_placeOpt_8),
    .f({_al_u1213_o,open_n3418}),
    .q({open_n3422,\picorv32_core/instr_bgeu }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(0*D*B*C*A)"),
    //.LUT1("(1*D*B*C*A)"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1214 (
    .a({_al_u1202_o,_al_u1202_o}),
    .b({_al_u1209_o,_al_u1209_o}),
    .c({_al_u1207_o,_al_u1207_o}),
    .d({_al_u1211_o,_al_u1211_o}),
    .mi({open_n3435,\picorv32_core/instr_beq }),
    .fx({open_n3440,_al_u1214_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(C*~(D*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b1010000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1216|picorv32_core/instr_bne_reg  (
    .a({\picorv32_core/alu_eq_lutinv ,\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .b({open_n3443,\picorv32_core/mem_rdata_q [12]}),
    .c({_al_u1215_o,\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_bne ,\picorv32_core/mem_rdata_q [14]}),
    .sr(resetn_placeOpt_8),
    .f({_al_u1216_o,open_n3456}),
    .q({open_n3460,\picorv32_core/instr_bne }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*~(B*~(A*~C)))"),
    //.LUTF1("B*C*~A*D+B*C*A*D"),
    //.LUTG0("(1*~D*~(B*~(A*~C)))"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000111011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1217|picorv32_core/mem_do_rinst_reg  (
    .a({open_n3461,\picorv32_core/n664_lutinv_placeOpt_7 }),
    .b({\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ,_al_u1552_o}),
    .c({\picorv32_core/n666_lutinv ,_al_u1555_o}),
    .clk(clk_pad),
    .d({resetn_placeOpt_17,_al_u1546_o}),
    .e({_al_u1216_o,resetn_placeOpt_17}),
    .sr(\picorv32_core/n728 ),
    .f({\picorv32_core/n728 ,open_n3477}),
    .q({open_n3481,\picorv32_core/mem_do_rinst }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D*~(~C*~B))"),
    //.LUT1("(A*~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))"),
    .INIT_LUT0(16'b0000000001010100),
    .INIT_LUT1(16'b0010000010101000),
    .MODE("LOGIC"))
    \_al_u1218|_al_u1219  (
    .a({_al_u1065_o,\uart/uart_status_rxd [3]}),
    .b({\uart/uart_status_rxd [0],\uart/n51_lutinv }),
    .c({rxd_pad,_al_u1065_o}),
    .d({\uart/mux37_b0_sel_is_3_o ,_al_u1218_o}),
    .f({_al_u1218_o,_al_u1219_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    .INIT_LUT0(16'b0011000000111111),
    .INIT_LUT1(16'b1111101000001010),
    .MODE("LOGIC"))
    \_al_u1220|_al_u1229  (
    .a({\uart/n49 [3],open_n3502}),
    .b({open_n3503,\uart/uart_smp_rx [0]}),
    .c({rxd_pad,rxd_pad}),
    .d({\uart/uart_smp_rx [3],\uart/n49 [0]}),
    .f({\uart/n50 [3],_al_u1229_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~(D*B)*~(~C*~A))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0011001011111010),
    .MODE("LOGIC"))
    \_al_u1221|_al_u1070  (
    .a({_al_u1068_o,open_n3524}),
    .b({\uart/n51_lutinv ,open_n3525}),
    .c({\uart/uart_smp_rx [3],\uart/uart_status_rxd [3]}),
    .d({_al_u1065_o,_al_u1065_o}),
    .f({_al_u1221_o,_al_u1070_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("B*~D*~C*~A+B*D*~C*~A+B*~D*C*~A+B*~D*~C*A+B*D*~C*A+B*~D*C*A"),
    //.LUTF1("A*~C*~B*~D+A*~C*B*~D+A*~C*~B*D+A*~C*B*D"),
    //.LUTG0("~B*~D*~C*~A+B*~D*~C*~A+~B*D*~C*~A+B*D*~C*~A+~B*~D*C*~A+B*~D*C*~A+~B*~D*~C*A+B*~D*~C*A+~B*D*~C*A+B*D*~C*A+~B*~D*C*A+B*~D*C*A"),
    //.LUTG1("A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b0000101000001010),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b1111101011111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1223|_al_u1224  (
    .a({\uart/n49 [2],open_n3546}),
    .b({open_n3547,_al_u1068_o}),
    .c({rxd_pad,_al_u1065_o}),
    .d({open_n3550,\uart/n51_lutinv }),
    .e({\uart/uart_smp_rx [2],\uart/uart_smp_rx [2]}),
    .f({\uart/n50 [2],_al_u1224_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A"),
    //.LUTF1("0"),
    //.LUTG0("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A"),
    //.LUTG1("~A*D*~C*~B+~A*D*~C*B"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000010100000101),
    .INIT_LUTG1(16'b0000010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1230|_al_u1068  (
    .a({\uart/uart_status_rxd [0],\uart/uart_status_rxd [0]}),
    .c({\uart/uart_status_rxd [2],\uart/uart_status_rxd [2]}),
    .d({\uart/uart_status_rxd [1],open_n3575}),
    .e({_al_u1229_o,\uart/uart_status_rxd [1]}),
    .f({_al_u1230_o,_al_u1068_o}));
  // ../src/uart.v(263)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(C)*~(D)*~((~0*B))+A*C*~(D)*~((~0*B))+A*C*D*~((~0*B))+A*~(C)*~(D)*(~0*B)+~(A)*C*~(D)*(~0*B)+A*C*~(D)*(~0*B)+~(A)*~(C)*D*(~0*B)+A*~(C)*D*(~0*B)+~(A)*C*D*(~0*B)+A*C*D*(~0*B))"),
    //.LUTF1("0"),
    //.LUTG0("(A*~(C)*~(D)*~((~1*B))+A*C*~(D)*~((~1*B))+A*C*D*~((~1*B))+A*~(C)*~(D)*(~1*B)+~(A)*C*~(D)*(~1*B)+A*C*~(D)*(~1*B)+~(A)*~(C)*D*(~1*B)+A*~(C)*D*(~1*B)+~(A)*C*D*(~1*B)+A*C*D*(~1*B))"),
    //.LUTG1("~A*D*~B*~C+~A*D*B*~C+~A*~D*~B*C+~A*D*~B*C+~A*~D*B*C+~A*D*B*C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110110011101010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010000010101010),
    .INIT_LUTG1(16'b0101010101010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1231|uart/reg9_b0  (
    .a({_al_u1230_o,_al_u1231_o}),
    .b({open_n3596,_al_u1232_o}),
    .c({_al_u1068_o,\uart/mux42_b0/B1_1 }),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({\uart/uart_smp_rx [0],_al_u1065_o}),
    .e({\uart/uart_status_rxd [3],\uart/uart_status_rxd [3]}),
    .sr(resetn_placeOpt_9),
    .f({_al_u1231_o,open_n3611}),
    .q({open_n3615,\uart/uart_smp_rx [0]}));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+~(A)*B*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+A*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0)"),
    //.LUT1("(~(C)*~(B)*~(A)*~(D)*~(1)+C*~(B)*~(A)*~(D)*~(1)+~(C)*B*~(A)*~(D)*~(1)+C*B*~(A)*~(D)*~(1)+~(C)*~(B)*A*~(D)*~(1)+C*~(B)*A*~(D)*~(1)+~(C)*B*A*~(D)*~(1)+C*B*A*~(D)*~(1)+~(C)*~(B)*~(A)*D*~(1)+C*~(B)*~(A)*D*~(1)+~(C)*~(B)*A*D*~(1)+~(C)*~(B)*~(A)*~(D)*1+C*~(B)*~(A)*~(D)*1+~(C)*B*~(A)*~(D)*1+C*B*~(A)*~(D)*1+~(C)*~(B)*A*~(D)*1+C*~(B)*A*~(D)*1+C*B*A*~(D)*1+~(C)*~(B)*~(A)*D*1+C*~(B)*~(A)*D*1+~(C)*~(B)*A*D*1)"),
    .INIT_LUT0(16'b0001001111111111),
    .INIT_LUT1(16'b0001001111110111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1232 (
    .a({\uart/uart_status_rxd [0],\uart/mux37_b0_sel_is_3_o }),
    .b({_al_u1229_o,_al_u1229_o}),
    .c({\uart/mux37_b0_sel_is_3_o ,\uart/uart_status_rxd [0]}),
    .d({rxd_pad,rxd_pad}),
    .mi({open_n3628,_al_u1065_o}),
    .fx({open_n3633,_al_u1232_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTF1("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG0("0"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*~C*B*D+A*~C*B*D"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1233|_al_u1065  (
    .a({_al_u1229_o,open_n3636}),
    .c({rxd_pad,\uart/uart_status_rxd [2]}),
    .e({\uart/n51_lutinv ,\uart/uart_status_rxd [1]}),
    .f({\uart/mux42_b0/B1_1 ,_al_u1065_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~A)"),
    //.LUT1("(D*C*~B*~A)"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0001000000000000),
    .MODE("LOGIC"))
    \_al_u1235|_al_u1238  (
    .a({\uart/n57 [4],\uart/n57 [4]}),
    .b({\uart/n57 [3],\uart/n57 [3]}),
    .c({\uart/n57 [2],\uart/n57 [2]}),
    .d({\uart/n51_lutinv ,\uart/n51_lutinv }),
    .f({_al_u1235_o,_al_u1238_o}));
  // ../src/uart.v(263)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(D)*~((~C*B*A))+0*D*~((~C*B*A))+~(0)*D*(~C*B*A)+0*D*(~C*B*A))"),
    //.LUTF1("~(0*~(C)*~((~D*~B*A))+0*C*~((~D*~B*A))+~(0)*C*(~D*~B*A)+0*C*(~D*~B*A))"),
    //.LUTG0("~(1*~(D)*~((~C*B*A))+1*D*~((~C*B*A))+~(1)*D*(~C*B*A)+1*D*(~C*B*A))"),
    //.LUTG1("~(1*~(C)*~((~D*~B*A))+1*C*~((~D*~B*A))+~(1)*C*(~D*~B*A)+1*C*(~D*~B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011111111111),
    .INIT_LUTF1(16'b1111111111011111),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1247|uart/reg6_b2  (
    .a({_al_u1238_o,_al_u1238_o}),
    .b({\uart/n57 [1],\uart/n57 [1]}),
    .c({_al_u1086_o,\uart/n57 [0]}),
    .ce(\uart/mux51_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\uart/n57 [0],_al_u1086_o}),
    .e({\uart/uart_idr_t [0],\uart/uart_idr_t [2]}),
    .mi({open_n3684,\uart/uart_idr_t [2]}),
    .sr(resetn_placeOpt_9),
    .f({_al_u1247_o,_al_u1243_o}),
    .q({open_n3699,\uart/uart_idr [2]}));  // ../src/uart.v(263)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~B*~A*~C*D)"),
    //.LUTF1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B"),
    //.LUTG0("(~1*~B*~A*~C*D)"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0011001100110011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1253|_al_u1123  (
    .a({open_n3700,\picorv32_core/n30 [17]}),
    .b({\picorv32_core/n30 [16],\picorv32_core/n30 [16]}),
    .c({open_n3701,\picorv32_core/n30 [18]}),
    .d({open_n3704,_al_u1122_o}),
    .e({\picorv32_core/n30 [14],\picorv32_core/n30 [14]}),
    .f({_al_u1253_o,_al_u1123_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~C*~B*A*D)"),
    //.LUTF1("(~0*~(~B*~A*D*C))"),
    //.LUTG0("(1*~C*~B*A*D)"),
    //.LUTG1("(~1*~(~B*~A*D*C))"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1110111111111111),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1254|_al_u1255  (
    .a({\picorv32_core/n30 [18],_al_u1175_o}),
    .b({\picorv32_core/n30 [17],_al_u1254_o}),
    .c({_al_u1253_o,_al_u1119_o}),
    .d({_al_u1122_o,_al_u1168_o}),
    .e({_al_u1121_o,_al_u1172_o}),
    .f({_al_u1254_o,uart_sel_lutinv}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~A*~C*B*D)"),
    //.LUTF1("(~0*~(~D*~C*B*A))"),
    //.LUTG0("(1*~A*~C*B*D)"),
    //.LUTG1("(~1*~(~D*~C*B*A))"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111111111110111),
    .INIT_LUTG0(16'b0000010000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1254|_al_u1255_placeOpt_1  (
    .a({_al_u1253_o,_al_u1119_o}),
    .b({_al_u1122_o,_al_u1175_o}),
    .c({\picorv32_core/n30 [18],_al_u1254_o}),
    .d({\picorv32_core/n30 [17],_al_u1168_o}),
    .e({_al_u1121_o,_al_u1172_o}),
    .f({open_n3764,uart_sel_lutinv_placeOpt_1}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~A*~B*C*D)"),
    //.LUTF1("(~0*~(~D*~C*B*A))"),
    //.LUTG0("(1*~A*~B*C*D)"),
    //.LUTG1("(~1*~(~D*~C*B*A))"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111111111110111),
    .INIT_LUTG0(16'b0001000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1254|_al_u1255_placeOpt_2  (
    .a({_al_u1253_o,_al_u1119_o}),
    .b({_al_u1122_o,_al_u1254_o}),
    .c({\picorv32_core/n30 [18],_al_u1175_o}),
    .d({\picorv32_core/n30 [17],_al_u1168_o}),
    .e({_al_u1121_o,_al_u1172_o}),
    .f({open_n3787,uart_sel_lutinv_placeOpt_2}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~A*~B*C*D)"),
    //.LUTF1("(~0*~(~C*~D*A*B))"),
    //.LUTG0("(1*~A*~B*C*D)"),
    //.LUTG1("(~1*~(~C*~D*A*B))"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111111111110111),
    .INIT_LUTG0(16'b0001000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1254|_al_u1255_placeOpt_3  (
    .a({_al_u1122_o,_al_u1119_o}),
    .b({_al_u1253_o,_al_u1254_o}),
    .c({\picorv32_core/n30 [17],_al_u1175_o}),
    .d({\picorv32_core/n30 [18],_al_u1168_o}),
    .e({_al_u1121_o,_al_u1172_o}),
    .f({open_n3810,uart_sel_lutinv_placeOpt_3}));
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~(A*~((B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D))*~(C)+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*~(C)+~(A)*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C)"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~(A*~((B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D))*~(C)+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*~(C)+~(A)*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111010100110101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0000010100110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1257|uart/reg0_b22  (
    .a({\picorv32_core/mem_rdata_q [22],\picorv32_core/pcpi_rs1$3$ }),
    .b({memory_out[22],\picorv32_core/n30 [1]}),
    .c({\picorv32_core/mem_xfer_placeOpt_4 ,_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_2,mem_la_addr[2]}),
    .e({uart_do[22],\uart/uart_bsrr [22]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1257_o,open_n3830}),
    .q({open_n3834,uart_do[22]}));  // ../src/uart.v(102)
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~0*~((~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))*~(A)+~0*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)*~(A)+~(~0)*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)*A+~0*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)*A)"),
    //.LUTF1("~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("~(~1*~((~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))*~(A)+~1*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)*~(A)+~(~1)*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)*A+~1*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)*A)"),
    //.LUTG1("D*B*~C*~A+~D*~B*C*~A+~D*B*C*~A+D*B*C*~A+D*B*~C*A+~D*~B*C*A+~D*B*C*A+D*B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000010101000),
    .INIT_LUTF1(16'b1010101010101010),
    .INIT_LUTG0(16'b0111010111111101),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1260|picorv32_core/reg0_b5  (
    .a({\picorv32_core/mem_rdata_q [5],\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({uart_do[5],_al_u1088_o}),
    .c({memory_out[5],\picorv32_core/mem_rdata_latched_noshuffle [5]}),
    .ce(\picorv32_core/mem_xfer ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_2,_al_u1261_o}),
    .e({\picorv32_core/mem_xfer ,\picorv32_core/mem_16bit_buffer [5]}),
    .f({\picorv32_core/mem_rdata_latched_noshuffle [5],\picorv32_core/mem_rdata_latched [5]}),
    .q({open_n3853,\picorv32_core/mem_rdata_q [5]}));  // ../src/picorv32.v(508)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~(A*~((B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D))*~(C)+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*~(C)+~(A)*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C)"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~(A*~((B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D))*~(C)+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*~(C)+~(A)*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111010100110101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0000010100110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1261|uart/reg0_b21  (
    .a({\picorv32_core/mem_rdata_q [21],\picorv32_core/pcpi_rs1$3$ }),
    .b({memory_out[21],\picorv32_core/n30 [1]}),
    .c({\picorv32_core/mem_xfer_placeOpt_4 ,_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_2,mem_la_addr[2]}),
    .e({uart_do[21],\uart/uart_bsrr [21]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1261_o,open_n3868}),
    .q({open_n3872,uart_do[21]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*C*~(A)*~(0)+~(B)*~(D)*~(C)*A*~(0)+~(B)*~(D)*C*A*~(0)+B*~(D)*C*A*~(0)+~(B)*D*~(C)*~(A)*0+B*~(D)*C*~(A)*0+~(B)*D*C*~(A)*0+~(B)*~(D)*~(C)*A*0+~(B)*D*~(C)*A*0+~(B)*~(D)*C*A*0+B*~(D)*C*A*0+~(B)*D*C*A*0)"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(B*~(D)*C*~(A)*~(1)+~(B)*~(D)*~(C)*A*~(1)+~(B)*~(D)*C*A*~(1)+B*~(D)*C*A*~(1)+~(B)*D*~(C)*~(A)*1+B*~(D)*C*~(A)*1+~(B)*D*C*~(A)*1+~(B)*~(D)*~(C)*A*1+~(B)*D*~(C)*A*1+~(B)*~(D)*C*A*1+B*~(D)*C*A*1+~(B)*D*C*A*1)"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011100010),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0011001111100010),
    .INIT_LUTG1(16'b1010101011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1263|uart/reg0_b4  (
    .a({uart_do[4],\uart/uart_odr [4]}),
    .b({\picorv32_core/mem_rdata_q [4],mem_la_addr[3]}),
    .c({memory_out[4],\uart/uart_bsrr [4]}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_xfer_placeOpt_1 ,mem_la_addr[2]}),
    .e({uart_sel_lutinv_placeOpt_1,\uart/uart_idr [4]}),
    .sr(resetn_placeOpt_13),
    .f({\picorv32_core/mem_rdata_latched_noshuffle [4],open_n3887}),
    .q({open_n3891,uart_do[4]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~D*~C*~B*~A+D*~C*~B*~A+~D*C*~B*~A+D*C*~B*~A+~D*~C*B*~A+D*~C*B*~A+~D*C*B*~A+D*C*B*~A"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~D*~C*~B*~A+D*~C*~B*~A+D*C*~B*~A+~D*~C*B*~A+~D*~C*~B*A+D*~C*~B*A+D*C*~B*A+~D*~C*B*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0011001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1264|uart/reg0_b20  (
    .a({\picorv32_core/mem_rdata_q [20],\picorv32_core/pcpi_rs1$3$ }),
    .b({uart_do[20],\picorv32_core/n30 [1]}),
    .c({memory_out[20],_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_2,mem_la_addr[2]}),
    .e({\picorv32_core/mem_xfer_placeOpt_1 ,\uart/uart_bsrr [20]}),
    .sr(resetn_placeOpt_13),
    .f({_al_u1264_o,open_n3906}),
    .q({open_n3910,uart_do[20]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*D*C*~B+A*D*C*~B+~A*~D*~C*B+A*~D*~C*B"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+~A*D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+~A*D*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0011001100001111),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0101010100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1266|uart/reg0_b19  (
    .a({uart_do[19],\picorv32_core/pcpi_rs1$3$ }),
    .b({memory_out[19],\picorv32_core/n30 [1]}),
    .c({\picorv32_core/mem_rdata_q [19],_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_xfer_placeOpt_1 ,mem_la_addr[2]}),
    .e({uart_sel_lutinv_placeOpt_1,\uart/uart_bsrr [19]}),
    .sr(resetn_placeOpt_13),
    .f({_al_u1266_o,open_n3925}),
    .q({open_n3929,uart_do[19]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*C*~(A)*~(0)+~(D)*~(B)*~(C)*A*~(0)+~(D)*~(B)*C*A*~(0)+D*~(B)*C*A*~(0)+~(D)*B*~(C)*~(A)*0+D*~(B)*C*~(A)*0+~(D)*B*C*~(A)*0+~(D)*~(B)*~(C)*A*0+~(D)*B*~(C)*A*0+~(D)*~(B)*C*A*0+D*~(B)*C*A*0+~(D)*B*C*A*0)"),
    //.LUTF1("(A*~((B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D))*~(C)+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*~(C)+~(A)*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C)"),
    //.LUTG0("(D*~(B)*C*~(A)*~(1)+~(D)*~(B)*~(C)*A*~(1)+~(D)*~(B)*C*A*~(1)+D*~(B)*C*A*~(1)+~(D)*B*~(C)*~(A)*1+D*~(B)*C*~(A)*1+~(D)*B*C*~(A)*1+~(D)*~(B)*~(C)*A*1+~(D)*B*~(C)*A*1+~(D)*~(B)*C*A*1+D*~(B)*C*A*1+~(D)*B*C*A*1)"),
    //.LUTG1("(A*~((B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D))*~(C)+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*~(C)+~(A)*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000000100010),
    .INIT_LUTF1(16'b0000101011001010),
    .INIT_LUTG0(16'b0011000011101110),
    .INIT_LUTG1(16'b1111101011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1267|uart/reg0_b3  (
    .a({\picorv32_core/mem_rdata_q [3],\uart/uart_odr [3]}),
    .b({memory_out[3],mem_la_addr[2]}),
    .c({\picorv32_core/mem_xfer_placeOpt_5 ,\uart/uart_bsrr [3]}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_3,mem_la_addr[3]}),
    .e({uart_do[3],\uart/uart_idr [3]}),
    .sr(resetn_placeOpt_15),
    .f({\picorv32_core/mem_rdata_latched_noshuffle [3],open_n3944}),
    .q({open_n3948,uart_do[3]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*~C*B+A*D*~C*B"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+~A*D*~C*B+~A*D*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0101010100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1270|uart/reg0_b18  (
    .a({uart_do[18],\picorv32_core/pcpi_rs1$3$ }),
    .b({\picorv32_core/mem_rdata_q [18],\picorv32_core/n30 [1]}),
    .c({memory_out[18],_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_xfer_placeOpt_1 ,mem_la_addr[2]}),
    .e({uart_sel_lutinv_placeOpt_1,\uart/uart_bsrr [18]}),
    .sr(resetn_placeOpt_13),
    .f({_al_u1270_o,open_n3963}),
    .q({open_n3967,uart_do[18]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*~B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0011001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1272|uart/reg0_b28  (
    .a({\picorv32_core/mem_rdata_q [28],\picorv32_core/pcpi_rs1$3$ }),
    .b({uart_do[28],\picorv32_core/n30 [1]}),
    .c({memory_out[28],_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_2,mem_la_addr[2]}),
    .e({\picorv32_core/mem_xfer_placeOpt_1 ,\uart/uart_bsrr [28]}),
    .sr(resetn_placeOpt_13),
    .f({_al_u1272_o,open_n3982}),
    .q({open_n3986,uart_do[28]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~C*~D*~A*~B+C*~D*~A*~B+~C*D*~A*~B+~C*~D*A*~B+C*~D*A*~B+~C*D*A*~B+~C*D*~A*B+~C*D*A*B"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~C*~D*~A*~B+C*~D*~A*~B+~C*D*~A*~B+C*D*~A*~B+~C*~D*A*~B+C*~D*A*~B+~C*D*~A*B+C*D*~A*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0101010100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1273|uart/reg0_b12  (
    .a({uart_do[12],\picorv32_core/pcpi_rs1$3$ }),
    .b({\picorv32_core/mem_rdata_q [12],\picorv32_core/n30 [1]}),
    .c({memory_out[12],_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_xfer_placeOpt_1 ,mem_la_addr[2]}),
    .e({uart_sel_lutinv_placeOpt_1,\uart/uart_bsrr [12]}),
    .sr(resetn_placeOpt_13),
    .f({_al_u1273_o,open_n4001}),
    .q({open_n4005,uart_do[12]}));  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~((B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D))*~(C)+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*~(C)+~(A)*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C)"),
    //.LUT1("(B*~((A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D))*~(C)+B*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)*~(C)+~(B)*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)*C+B*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)*C)"),
    .INIT_LUT0(16'b0000101011001010),
    .INIT_LUT1(16'b1111110010101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1275 (
    .a({memory_out[1],\picorv32_core/mem_rdata_q [1]}),
    .b({\picorv32_core/mem_rdata_q [1],memory_out[1]}),
    .c({\picorv32_core/mem_xfer_placeOpt_5 ,\picorv32_core/mem_xfer_placeOpt_5 }),
    .d({uart_sel_lutinv_placeOpt_3,uart_sel_lutinv_placeOpt_3}),
    .mi({open_n4018,uart_do[1]}),
    .fx({open_n4023,\picorv32_core/mem_rdata_latched_noshuffle [1]}));
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~(A*~((B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D))*~(C)+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*~(C)+~(A)*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C)"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~(A*~((B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D))*~(C)+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*~(C)+~(A)*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111010100110101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0000010100110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1276|uart/reg0_b17  (
    .a({\picorv32_core/mem_rdata_q [17],\picorv32_core/pcpi_rs1$3$ }),
    .b({memory_out[17],\picorv32_core/n30 [1]}),
    .c({\picorv32_core/mem_xfer_placeOpt_5 ,_al_u700_o_placeOpt_2}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_3,mem_la_addr[2]}),
    .e({uart_do[17],\uart/uart_bsrr [17]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1276_o,open_n4040}),
    .q({open_n4044,uart_do[17]}));  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*A*~D*~(~0*~C))"),
    //.LUTF1("~C*~B*~D*~A+C*~B*~D*~A+~C*B*~D*~A+C*B*~D*~A+~C*~B*D*~A+C*~B*D*~A+~C*B*~D*A+C*B*~D*A"),
    //.LUTG0("(~B*A*~D*~(~1*~C))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b0001000111011101),
    .INIT_LUTG0(16'b0000000000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1278|_al_u1279  (
    .a({\picorv32_core/n30 [6],_al_u1278_o}),
    .b({_al_u700_o,\eq2/or_xor_i0$1$_i1$1$_o_o_lutinv }),
    .c({open_n4045,_al_u1123_o}),
    .d({\picorv32_core/pcpi_rs1$8$ ,_al_u1119_o}),
    .e({mem_la_addr[7],_al_u1121_o}),
    .f({_al_u1278_o,_al_u1279_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(0)*~((A*D*C))+B*0*~((A*D*C))+~(B)*0*(A*D*C)+B*0*(A*D*C))"),
    //.LUTF1("(B*~(0)*~((A*D*C))+B*0*~((A*D*C))+~(B)*0*(A*D*C)+B*0*(A*D*C))"),
    //.LUTG0("(B*~(1)*~((A*D*C))+B*1*~((A*D*C))+~(B)*1*(A*D*C)+B*1*(A*D*C))"),
    //.LUTG1("(B*~(1)*~((A*D*C))+B*1*~((A*D*C))+~(B)*1*(A*D*C)+B*1*(A*D*C))"),
    .INIT_LUTF0(16'b0100110011001100),
    .INIT_LUTF1(16'b0100110011001100),
    .INIT_LUTG0(16'b1110110011001100),
    .INIT_LUTG1(16'b1110110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1280|_al_u1525  (
    .a({_al_u1175_o,_al_u1175_o}),
    .b({memory_out[1],memory_out[27]}),
    .c({_al_u1279_o,_al_u1279_o}),
    .d({_al_u1168_o,_al_u1168_o}),
    .e({uart_do[1],uart_do[27]}),
    .f({mem_rdata[1],mem_rdata[27]}));
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0011001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1282|uart/reg0_b16  (
    .a({\picorv32_core/mem_rdata_q [16],\picorv32_core/pcpi_rs1$3$ }),
    .b({uart_do[16],\picorv32_core/n30 [1]}),
    .c({memory_out[16],_al_u700_o_placeOpt_2}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_3,mem_la_addr[2]}),
    .e({\picorv32_core/mem_xfer_placeOpt_5 ,\uart/uart_bsrr [16]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1282_o,open_n4104}),
    .q({open_n4108,uart_do[16]}));  // ../src/uart.v(102)
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*D*(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A))"),
    //.LUTF1("~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("~(~B*D*(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A))"),
    //.LUTG1("D*B*~C*~A+~D*~B*C*~A+~D*B*C*~A+D*B*C*~A+D*B*~C*A+~D*~B*C*A+~D*B*C*A+D*B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110111111111111),
    .INIT_LUTF1(16'b1010101010101010),
    .INIT_LUTG0(16'b1100110111111111),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1283|picorv32_core/prefetched_high_word_reg  (
    .a({\picorv32_core/mem_rdata_q [0],uart_sel_lutinv_placeOpt_3}),
    .b({uart_do[0],\picorv32_core/mem_la_secondword }),
    .c({memory_out[0],memory_out[0]}),
    .ce(\picorv32_core/mux61_sel_is_5_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_3,mem_rdata[1]}),
    .e({\picorv32_core/mem_xfer_placeOpt_5 ,uart_do[0]}),
    .sr(\picorv32_core/u179_sel_is_0_o ),
    .f({\picorv32_core/mem_rdata_latched_noshuffle [0],\picorv32_core/n131 }),
    .q({open_n4126,\picorv32_core/prefetched_high_word }));  // ../src/picorv32.v(605)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*D)"),
    //.LUTF1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+A*~D*C*B"),
    //.LUTG0("~(~C*D)"),
    //.LUTG1("A*~D*~C*~B+A*D*~C*~B+A*~D*C*~B+A*~D*~C*B+A*D*~C*B+A*~D*C*B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111111),
    .INIT_LUTF1(16'b0000111111111111),
    .INIT_LUTG0(16'b1111000011111111),
    .INIT_LUTG1(16'b0000101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1285|picorv32_core/is_lui_auipc_jal_reg  (
    .a({_al_u1151_o,open_n4127}),
    .c({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .clk(clk_pad),
    .d({\picorv32_core/sel39_b0_sel_is_3_o ,_al_u665_o}),
    .e({\picorv32_core/latched_branch ,open_n4131}),
    .f({_al_u1285_o,\picorv32_core/n472 }),
    .q({open_n4150,\picorv32_core/is_lui_auipc_jal }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~B*~A*~D*~C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1288|picorv32_core/reg19_b32  (
    .a({\picorv32_core/instr_rdinstr ,\picorv32_core/instr_rdcycle }),
    .b({\picorv32_core/instr_rdinstrh ,\picorv32_core/instr_rdinstrh }),
    .c({\picorv32_core/instr_rdcycle ,\picorv32_core/count_cycle [0]}),
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_rdcycleh ,\picorv32_core/count_instr [32]}),
    .mi({open_n4161,\picorv32_core/n503 [32]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1288_o,_al_u1902_o}),
    .q({open_n4165,\picorv32_core/count_instr [32]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("(~A*~(~0*~D*~C*~B))"),
    //.LUTG0("A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG1("(~A*~(~1*~D*~C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110111011101110),
    .INIT_LUTF1(16'b0101010101010100),
    .INIT_LUTG0(16'b1010111010101110),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1290|picorv32_core/latched_store_reg  (
    .a({_al_u1151_o,_al_u1290_o}),
    .b({\picorv32_core/sel40_b6/B5 ,\picorv32_core/n666_lutinv }),
    .c({\picorv32_core/n669_lutinv ,\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .clk(clk_pad),
    .d({\picorv32_core/n667_lutinv ,open_n4167}),
    .e({\picorv32_core/latched_store ,_al_u1216_o}),
    .sr(resetn_placeOpt_10),
    .f({_al_u1290_o,open_n4182}),
    .q({open_n4186,\picorv32_core/latched_store }));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("(~D*~(0*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)))"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("(~D*~(1*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)))"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b0000000000011011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1293|_al_u1292  (
    .a({\picorv32_core/instr_sub ,_al_u826_o}),
    .b({\picorv32_core/n434 [0],_al_u827_o}),
    .c({\picorv32_core/n433 [0],_al_u828_o}),
    .d({_al_u1292_o,\picorv32_core/pcpi_rs1$0$ }),
    .e({\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub ,mem_la_wdata[0]}),
    .f({_al_u1293_o,_al_u1292_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*B)"),
    //.LUTF1("~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    //.LUTG0("(D*B)"),
    //.LUTG1("~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    .INIT_LUTF0(16'b1100110000000000),
    .INIT_LUTF1(16'b1100110011001100),
    .INIT_LUTG0(16'b1100110000000000),
    .INIT_LUTG1(16'b1100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1295|_al_u1115  (
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mem_xfer }),
    .c({_al_u1276_o,open_n4211}),
    .d({open_n4214,_al_u1088_o}),
    .e({_al_u1088_o,open_n4215}),
    .f({_al_u1295_o,\picorv32_core/mem_la_firstword_xfer }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~C*~B)"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"))
    \_al_u1296|_al_u1638  (
    .a({open_n4236,\picorv32_core/mem_16bit_buffer [13]}),
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .c({\picorv32_core/mem_16bit_buffer [1],open_n4237}),
    .f({_al_u1296_o,_al_u1638_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*B*A)"),
    //.LUT1("(~A*~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1298|picorv32_core/instr_bge_reg  (
    .a({\picorv32_core/instr_xori ,\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .b({\picorv32_core/instr_bge ,\picorv32_core/mem_rdata_q [12]}),
    .c({\picorv32_core/instr_xor ,\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_beq ,\picorv32_core/mem_rdata_q [14]}),
    .sr(resetn_placeOpt_8),
    .f({_al_u1298_o,open_n4272}),
    .q({open_n4276,\picorv32_core/instr_bge }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("0"),
    //.LUTG0("D*~B*~C*~A+D*~B*~C*A"),
    //.LUTG1("~C*~D*~A*~B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1299|picorv32_core/instr_blt_reg  (
    .a({\picorv32_core/instr_blt ,open_n4277}),
    .b({\picorv32_core/instr_bltu ,\picorv32_core/mem_rdata_q [12]}),
    .c({\picorv32_core/instr_bne ,\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_bgeu ,\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .e({_al_u1298_o,\picorv32_core/mem_rdata_q [14]}),
    .sr(resetn_placeOpt_8),
    .f({_al_u1299_o,open_n4292}),
    .q({open_n4296,\picorv32_core/instr_blt }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~A*~D*~C*~B+~A*~D*~C*B"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000101),
    .INIT_LUTG0(16'b0000000000001010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1300|picorv32_core/instr_sh_reg  (
    .a({\picorv32_core/instr_sb ,\picorv32_core/is_sb_sh_sw }),
    .c({\picorv32_core/instr_lb ,\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sh ,\picorv32_core/mem_rdata_q [14]}),
    .e({\picorv32_core/instr_lh ,\picorv32_core/mem_rdata_q [12]}),
    .f({_al_u1300_o,open_n4314}),
    .q({open_n4318,\picorv32_core/instr_sh }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(~0*~B*~A*C*D)"),
    //.LUTG0("A*~B*~C*D+A*B*~C*D"),
    //.LUTG1("(~1*~B*~A*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0000101000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1301|picorv32_core/instr_srl_reg  (
    .a({\picorv32_core/instr_srl ,_al_u976_o}),
    .b({\picorv32_core/instr_srli ,open_n4319}),
    .c({_al_u1300_o,\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({_al_u1299_o,\picorv32_core/mem_rdata_q [14]}),
    .e({\picorv32_core/instr_sw ,\picorv32_core/mem_rdata_q [12]}),
    .sr(resetn_placeOpt_16),
    .f({_al_u1301_o,open_n4334}),
    .q({open_n4338,\picorv32_core/instr_srl }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*C*B*A)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~1*~D*C*B*A)"),
    //.LUTG1("(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1302|picorv32_core/instr_sll_reg  (
    .a({open_n4339,\picorv32_core/n304_lutinv }),
    .b({open_n4340,\picorv32_core/is_alu_reg_reg }),
    .c({\picorv32_core/instr_slli ,\picorv32_core/mem_rdata_q [12]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sll ,\picorv32_core/mem_rdata_q [13]}),
    .e({open_n4341,\picorv32_core/mem_rdata_q [14]}),
    .sr(resetn_placeOpt_17),
    .f({_al_u1302_o,open_n4356}),
    .q({open_n4360,\picorv32_core/instr_sll }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(~0*~A*C*B*D)"),
    //.LUTG0("~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG1("(~1*~A*C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0100000000000000),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1303|picorv32_core/instr_sra_reg  (
    .a({\picorv32_core/instr_sra ,open_n4361}),
    .b({_al_u828_o,\picorv32_core/is_alu_reg_reg }),
    .c({_al_u1302_o,open_n4362}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({_al_u827_o,open_n4363}),
    .e({\picorv32_core/instr_srai ,\picorv32_core/n345 }),
    .sr(resetn_placeOpt_8),
    .f({_al_u1303_o,open_n4378}),
    .q({open_n4382,\picorv32_core/instr_sra }));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~A*~C*~B*~D)"),
    //.LUTF1("(0*B*C*~D*A)"),
    //.LUTG0("(~1*~A*~C*~B*~D)"),
    //.LUTG1("(1*B*C*~D*A)"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1305|_al_u1304  (
    .a({_al_u1301_o,\picorv32_core/instr_sltiu }),
    .b({_al_u1304_o,\picorv32_core/instr_slt }),
    .c({_al_u1303_o,\picorv32_core/instr_slti }),
    .d({\picorv32_core/n165 ,\picorv32_core/n168 }),
    .e({_al_u1288_o,\picorv32_core/instr_sltu }),
    .f({\picorv32_core/n524 [7],_al_u1304_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("A*~C*~B*~D+A*C*~B*~D+A*~C*~B*D+A*C*~B*D"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTG1("A*~C*~B*~D+A*C*~B*~D+A*~C*~B*D+A*C*~B*D"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0010001000100010),
    .INIT_LUTG0(16'b0000111100001111),
    .INIT_LUTG1(16'b0010001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1306|_al_u1289  (
    .a({_al_u1288_o,open_n4405}),
    .b({\picorv32_core/is_slli_srli_srai ,open_n4406}),
    .c({open_n4407,_al_u1288_o}),
    .e({open_n4412,\picorv32_core/n664_lutinv_placeOpt_1 }),
    .f({_al_u1306_o,\picorv32_core/sel40_b6/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*~A)"),
    //.LUT1("(~1*~D*~C*~B*~A)"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1308 (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .mi({open_n4445,\picorv32_core/decoded_rs2 [4]}),
    .fx({open_n4450,_al_u1308_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0100010001010000),
    .MODE("LOGIC"))
    \_al_u1309|_al_u1327  (
    .a({_al_u1308_o,_al_u1308_o}),
    .b({\picorv32_core/cpuregs_p2/dram_do_i1_004 ,\picorv32_core/decoded_rs2 [4]}),
    .c({\picorv32_core/cpuregs_p2/dram_do_i0_004 ,\picorv32_core/cpuregs_p2/dram_do_i0_001 }),
    .d({\picorv32_core/decoded_rs2 [4],\picorv32_core/cpuregs_p2/dram_do_i1_001 }),
    .f({\picorv32_core/cpuregs_rs2 [4],\picorv32_core/cpuregs_rs2 [1]}));
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(C*~D)))"),
    //.LUT1("~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001010100010),
    .INIT_LUT1(16'b0101000001011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1310|picorv32_core/reg12_b4  (
    .a({\picorv32_core/cpuregs_rs2 [4],resetn_placeOpt_17}),
    .b({open_n4473,_al_u1315_o}),
    .c({\picorv32_core/n523_lutinv ,\picorv32_core/n664_lutinv_placeOpt_6 }),
    .clk(clk_pad),
    .d({\picorv32_core/decoded_rs2 [4],_al_u1310_o}),
    .f({_al_u1310_o,open_n4488}),
    .q({open_n4492,\picorv32_core/reg_sh [4]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~C*~B*A*D)"),
    //.LUT1("(~1*~D*~B*A*C)"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1311 (
    .a(2'b00),
    .b({\picorv32_core/cpu_state [5],\picorv32_core/cpu_state [5]}),
    .c({_al_u982_o,\picorv32_core/cpu_state [6]}),
    .d({\picorv32_core/cpu_state [6],_al_u982_o}),
    .mi({open_n4505,\picorv32_core/cpu_state [7]}),
    .fx({open_n4510,\picorv32_core/n665_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*A*~B*D+C*A*~B*D+~C*A*B*D+C*A*B*D"),
    //.LUTF1("(D*B)"),
    //.LUTG0("~C*A*B*~D+C*A*B*~D+~C*A*B*D+C*A*B*D"),
    //.LUTG1("(D*B)"),
    .INIT_LUTF0(16'b1010101000000000),
    .INIT_LUTF1(16'b1100110000000000),
    .INIT_LUTG0(16'b1000100010001000),
    .INIT_LUTG1(16'b1100110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1312|_al_u1355  (
    .a({open_n4513,\picorv32_core/n664_lutinv_placeOpt_6 }),
    .b({\picorv32_core/n665_lutinv ,\picorv32_core/cpuregs_rs2 [4]}),
    .d({\picorv32_core/cpuregs_rs2 [4],\picorv32_core/decoded_imm [4]}),
    .e({open_n4518,\picorv32_core/n523_lutinv }),
    .f({\picorv32_core/sel42_b4/B4 ,\picorv32_core/sel42_b4/B5 }));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A)"),
    //.LUTF1("(~0*~C*~D*~B*~A)"),
    //.LUTG0("(B*~A)"),
    //.LUTG1("(~1*~C*~D*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010001000100),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0100010001000100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1313|picorv32_core/reg12_b3  (
    .a({\picorv32_core/reg_sh [0],_al_u1320_o}),
    .b({\picorv32_core/reg_sh [1],resetn_placeOpt_17}),
    .c({\picorv32_core/reg_sh [3],open_n4539}),
    .clk(clk_pad),
    .d({\picorv32_core/reg_sh [2],open_n4541}),
    .e({\picorv32_core/reg_sh [4],open_n4542}),
    .f({_al_u1313_o,open_n4558}),
    .q({open_n4562,\picorv32_core/reg_sh [3]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(C*A*B)"),
    //.LUT1("(~A*B)"),
    .INIT_LUT0(16'b1000000010000000),
    .INIT_LUT1(16'b0100010001000100),
    .MODE("LOGIC"))
    \_al_u1314|_al_u1742  (
    .a({_al_u1313_o,_al_u1313_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .c({open_n4563,\picorv32_core/pcpi_rs1$29$ }),
    .f({\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv ,\picorv32_core/sel43_b29/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*D+~A*B*C*D"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0100010000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0101010100010001),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1318|_al_u1317  (
    .a({\picorv32_core/cpuregs_rs2 [3],_al_u1308_o}),
    .b({open_n4586,\picorv32_core/decoded_rs2 [4]}),
    .d({open_n4591,\picorv32_core/cpuregs_p2/dram_do_i1_003 }),
    .e({\picorv32_core/n665_lutinv ,\picorv32_core/cpuregs_p2/dram_do_i0_003 }),
    .f({\picorv32_core/sel42_b3/B4 ,\picorv32_core/cpuregs_rs2 [3]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(B*(0*~(D)*~(C)+0*D*~(C)+~(0)*D*C+0*D*C)))"),
    //.LUT1("(~A*~(B*(1*~(D)*~(C)+1*D*~(C)+~(1)*D*C+1*D*C)))"),
    .INIT_LUT0(16'b0001010101010101),
    .INIT_LUT1(16'b0001000101010001),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1319 (
    .a({\picorv32_core/sel42_b3/B4 ,\picorv32_core/sel42_b3/B4 }),
    .b({\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv ,\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv }),
    .c({\picorv32_core/n554 ,\picorv32_core/n554 }),
    .d({\picorv32_core/n559 [3],\picorv32_core/n559 [3]}),
    .mi({open_n4624,\picorv32_core/n564 [3]}),
    .fx({open_n4629,_al_u1319_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUT1("(B*~(C*(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .INIT_LUT0(16'b0100110011001100),
    .INIT_LUT1(16'b0000110010001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1320 (
    .a({\picorv32_core/n523_lutinv ,\picorv32_core/n523_lutinv }),
    .b({_al_u1319_o,_al_u1319_o}),
    .c({\picorv32_core/n664_lutinv_placeOpt_6 ,\picorv32_core/n664_lutinv_placeOpt_6 }),
    .d({\picorv32_core/cpuregs_rs2 [3],\picorv32_core/cpuregs_rs2 [3]}),
    .mi({open_n4644,\picorv32_core/decoded_rs2 [3]}),
    .fx({open_n4649,_al_u1320_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*D*~C+~A*~B*D*C"),
    //.LUTF1("(D*A)"),
    //.LUTG0("~A*B*~D*~C+~A*~B*D*~C+~A*B*D*~C+~A*B*~D*C+~A*~B*D*C+~A*B*D*C"),
    //.LUTG1("(D*A)"),
    .INIT_LUTF0(16'b0001000100000000),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b0101010101000100),
    .INIT_LUTG1(16'b1010101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1323|_al_u1322  (
    .a({\picorv32_core/n665_lutinv ,_al_u1308_o}),
    .b({open_n4652,\picorv32_core/decoded_rs2 [4]}),
    .d({\picorv32_core/cpuregs_rs2 [2],\picorv32_core/cpuregs_p2/dram_do_i0_002 }),
    .e({open_n4657,\picorv32_core/cpuregs_p2/dram_do_i1_002 }),
    .f({\picorv32_core/sel42_b2/B4 ,\picorv32_core/cpuregs_rs2 [2]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(B*(0*~(D)*~(C)+0*D*~(C)+~(0)*D*C+0*D*C)))"),
    //.LUT1("(~A*~(B*(1*~(D)*~(C)+1*D*~(C)+~(1)*D*C+1*D*C)))"),
    .INIT_LUT0(16'b0001010101010101),
    .INIT_LUT1(16'b0001000101010001),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1324 (
    .a({\picorv32_core/sel42_b2/B4 ,\picorv32_core/sel42_b2/B4 }),
    .b({\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv ,\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv }),
    .c({\picorv32_core/n554 ,\picorv32_core/n554 }),
    .d({\picorv32_core/n559 [2],\picorv32_core/n559 [2]}),
    .mi({open_n4690,\picorv32_core/n564 [2]}),
    .fx({open_n4695,_al_u1324_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(C*A)"),
    //.LUTG0("A*~D*C*~B+A*D*C*~B+~A*~D*~C*B+~A*D*~C*B+~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    //.LUTG1("(C*A)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010000010100000),
    .INIT_LUTG0(16'b1110010011100100),
    .INIT_LUTG1(16'b1010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1328|_al_u1397  (
    .a({\picorv32_core/n665_lutinv ,\picorv32_core/n523_lutinv }),
    .b({open_n4698,\picorv32_core/decoded_imm [1]}),
    .c({\picorv32_core/cpuregs_rs2 [1],\picorv32_core/cpuregs_rs2 [1]}),
    .e({open_n4703,\picorv32_core/n664_lutinv_placeOpt_3 }),
    .f({\picorv32_core/sel42_b1/B4 ,\picorv32_core/sel42_b1/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*D)"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1010101000000000),
    .MODE("LOGIC"))
    \_al_u1333|_al_u1332  (
    .a({\picorv32_core/cpuregs_rs2 [0],_al_u1308_o}),
    .b({open_n4724,\picorv32_core/decoded_rs2 [4]}),
    .c({open_n4725,\picorv32_core/cpuregs_p2/dram_do_i0_000 }),
    .d({\picorv32_core/n665_lutinv ,\picorv32_core/cpuregs_p2/dram_do_i1_000 }),
    .f({\picorv32_core/sel42_b0/B4 ,\picorv32_core/cpuregs_rs2 [0]}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~D)"),
    //.LUTF1("(~C*~(B*(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTG0("(A*~D)"),
    //.LUTG1("(~C*~(B*(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010101010),
    .INIT_LUTF1(16'b0000011100001111),
    .INIT_LUTG0(16'b0000000010101010),
    .INIT_LUTG1(16'b0000001100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1334|picorv32_core/reg12_b0  (
    .a({\picorv32_core/n554 ,resetn_placeOpt_17}),
    .b({\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv ,open_n4746}),
    .c({\picorv32_core/sel42_b0/B4 ,open_n4747}),
    .clk(clk_pad),
    .d({\picorv32_core/n559 [0],_al_u1335_o}),
    .e({\picorv32_core/n564 [0],open_n4749}),
    .f({_al_u1334_o,open_n4765}),
    .q({open_n4769,\picorv32_core/reg_sh [0]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUT1("(B*~(C*(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .INIT_LUT0(16'b0100110011001100),
    .INIT_LUT1(16'b0000110010001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1335 (
    .a({\picorv32_core/n523_lutinv ,\picorv32_core/n523_lutinv }),
    .b({_al_u1334_o,_al_u1334_o}),
    .c({\picorv32_core/n664_lutinv_placeOpt_6 ,\picorv32_core/n664_lutinv_placeOpt_6 }),
    .d({\picorv32_core/cpuregs_rs2 [0],\picorv32_core/cpuregs_rs2 [0]}),
    .mi({open_n4782,\picorv32_core/decoded_rs2 [0]}),
    .fx({open_n4787,_al_u1335_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTG0("0"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1337|_al_u2493  (
    .b({\picorv32_core/n664_lutinv_placeOpt_6 ,open_n4792}),
    .c({\picorv32_core/n665_lutinv ,open_n4793}),
    .e({\picorv32_core/n523_lutinv ,resetn_placeOpt_17}),
    .f({_al_u1337_o,\picorv32_core/n407 }));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*B*~D*A+C*B*~D*A+~C*B*D*A+C*B*D*A"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D"),
    //.LUTG0("~C*B*~D*A+C*B*~D*A+~C*~B*D*A+C*~B*D*A+~C*B*D*A+C*B*D*A"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b1010101010001000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1338|picorv32_core/reg22_b7  (
    .a({\picorv32_core/n663 ,resetn_placeOpt_8}),
    .b({open_n4818,\picorv32_core/n662 }),
    .clk(clk_pad),
    .d({\picorv32_core/n662 ,\picorv32_core/n664_lutinv_placeOpt_1 }),
    .e({\picorv32_core/n666_lutinv ,\picorv32_core/n524 [7]}),
    .sr(\picorv32_core/mux164_b0_sel_is_0_o ),
    .f({_al_u1338_o,open_n4836}),
    .q({open_n4840,\picorv32_core/cpu_state [7]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*~B)*~(D*C*~A))"),
    //.LUT1("(~(1*~D)*~(B*C*~A))"),
    .INIT_LUT0(16'b1010111111111111),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1340 (
    .a({\picorv32_core/n523_lutinv ,\picorv32_core/n523_lutinv }),
    .b({\picorv32_core/decoded_imm [9],_al_u1339_o}),
    .c({\picorv32_core/n664_lutinv_placeOpt_7 ,\picorv32_core/n664_lutinv_placeOpt_7 }),
    .d({_al_u1339_o,\picorv32_core/decoded_imm [9]}),
    .mi({open_n4853,\picorv32_core/pcpi_rs2$9$ }),
    .fx({open_n4858,_al_u1340_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~(D*~C))"),
    //.LUT1("(~A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101111101010101),
    .INIT_LUT1(16'b0100010001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1341|picorv32_core/reg26_b9  (
    .a({_al_u1308_o,_al_u1340_o}),
    .b({\picorv32_core/cpuregs_p2/dram_do_i1_009 ,open_n4861}),
    .c({\picorv32_core/cpuregs_p2/dram_do_i0_009 ,_al_u1337_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoded_rs2 [4],\picorv32_core/cpuregs_rs2 [9]}),
    .f({\picorv32_core/cpuregs_rs2 [9],open_n4875}),
    .q({open_n4879,\picorv32_core/pcpi_rs2$9$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0011001000000010),
    .MODE("LOGIC"))
    \_al_u1344|_al_u1424  (
    .a({\picorv32_core/cpuregs_p2/dram_do_i0_008 ,_al_u1308_o}),
    .b({_al_u1308_o,\picorv32_core/decoded_rs2 [4]}),
    .c({\picorv32_core/decoded_rs2 [4],\picorv32_core/cpuregs_p2/dram_do_i0_011 }),
    .d({\picorv32_core/cpuregs_p2/dram_do_i1_008 ,\picorv32_core/cpuregs_p2/dram_do_i1_011 }),
    .f({\picorv32_core/cpuregs_rs2 [8],\picorv32_core/cpuregs_rs2 [11]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*~B)*~(D*C*~A))"),
    //.LUT1("(~(1*~B)*~(A*C*~D))"),
    .INIT_LUT0(16'b1010111111111111),
    .INIT_LUT1(16'b1100110001001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1346 (
    .a({\picorv32_core/decoded_imm [7],\picorv32_core/n523_lutinv }),
    .b({_al_u1339_o,_al_u1339_o}),
    .c({\picorv32_core/n664_lutinv ,\picorv32_core/n664_lutinv }),
    .d({\picorv32_core/n523_lutinv ,\picorv32_core/decoded_imm [7]}),
    .mi({open_n4912,mem_la_wdata[7]}),
    .fx({open_n4917,_al_u1346_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("A*B*~C*~D+A*B*C*~D"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D+A*~B*~C*D+A*B*~C*D"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0000000010001000),
    .INIT_LUTG0(16'b0000101000001010),
    .INIT_LUTG1(16'b0000000011011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1347|picorv32_core/reg26_b7  (
    .a({\picorv32_core/decoded_rs2 [4],\picorv32_core/cpuregs_rs2 [7]}),
    .b({\picorv32_core/cpuregs_p2/dram_do_i1_007 ,open_n4920}),
    .c({open_n4921,_al_u1337_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1308_o,open_n4922}),
    .e({\picorv32_core/cpuregs_p2/dram_do_i0_007 ,_al_u1346_o}),
    .f({\picorv32_core/cpuregs_rs2 [7],open_n4938}),
    .q({open_n4942,mem_la_wdata[7]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0100010001010000),
    .MODE("LOGIC"))
    \_al_u1350|_al_u1421  (
    .a({_al_u1308_o,_al_u1308_o}),
    .b({\picorv32_core/cpuregs_p2/dram_do_i1_006 ,\picorv32_core/decoded_rs2 [4]}),
    .c({\picorv32_core/cpuregs_p2/dram_do_i0_006 ,\picorv32_core/cpuregs_p2/dram_do_i0_012 }),
    .d({\picorv32_core/decoded_rs2 [4],\picorv32_core/cpuregs_p2/dram_do_i1_012 }),
    .f({\picorv32_core/cpuregs_rs2 [6],\picorv32_core/cpuregs_rs2 [12]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~D*C+~A*B*D*C"),
    //.LUTF1("A*C*~D*~B+A*C*D*~B"),
    //.LUTG0("~A*~B*~D*~C+~A*~B*D*~C+~A*~B*~D*C+~A*B*~D*C+~A*~B*D*C+~A*B*D*C"),
    //.LUTG1("~A*~C*~D*~B+~A*C*~D*~B+A*C*~D*~B+~A*~C*D*~B+~A*C*D*~B+A*C*D*~B"),
    .INIT_LUTF0(16'b0100000001000000),
    .INIT_LUTF1(16'b0010000000100000),
    .INIT_LUTG0(16'b0101000101010001),
    .INIT_LUTG1(16'b0011000100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1353|_al_u1412  (
    .a({\picorv32_core/decoded_rs2 [4],_al_u1308_o}),
    .b({_al_u1308_o,\picorv32_core/decoded_rs2 [4]}),
    .c({\picorv32_core/cpuregs_p2/dram_do_i1_005 ,\picorv32_core/cpuregs_p2/dram_do_i1_015 }),
    .e({\picorv32_core/cpuregs_p2/dram_do_i0_005 ,\picorv32_core/cpuregs_p2/dram_do_i0_015 }),
    .f({\picorv32_core/cpuregs_rs2 [5],\picorv32_core/cpuregs_rs2 [15]}));
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D*~(A*~B))"),
    //.LUT1("(D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110010),
    .INIT_LUT1(16'b1110010000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1357|picorv32_core/reg26_b3  (
    .a({\picorv32_core/n523_lutinv ,mem_la_wdata[3]}),
    .b({\picorv32_core/decoded_imm [3],_al_u1339_o}),
    .c({\picorv32_core/cpuregs_rs2 [3],\picorv32_core/sel42_b3/B4 }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/n664_lutinv_placeOpt_6 ,\picorv32_core/sel42_b3/B5 }),
    .f({\picorv32_core/sel42_b3/B5 ,open_n5000}),
    .q({open_n5004,mem_la_wdata[3]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~A*D*~B+~C*~A*D*B"),
    //.LUTF1("~B*D*~C*A+B*D*~C*A"),
    //.LUTG0("~C*A*~D*~B+~C*~A*D*~B+~C*A*D*~B+~C*A*~D*B+~C*~A*D*B+~C*A*D*B"),
    //.LUTG1("~B*~D*~C*~A+B*~D*~C*~A+~B*~D*~C*A+B*~D*~C*A+~B*D*~C*A+B*D*~C*A"),
    .INIT_LUTF0(16'b0000010100000000),
    .INIT_LUTF1(16'b0000101000000000),
    .INIT_LUTG0(16'b0000111100001010),
    .INIT_LUTG1(16'b0000101000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1360|_al_u1406  (
    .a({\picorv32_core/cpuregs_p2/dram_do_i1_031 ,\picorv32_core/decoded_rs2 [4]}),
    .c({_al_u1308_o,_al_u1308_o}),
    .d({\picorv32_core/decoded_rs2 [4],\picorv32_core/cpuregs_p2/dram_do_i0_017 }),
    .e({\picorv32_core/cpuregs_p2/dram_do_i0_031 ,\picorv32_core/cpuregs_p2/dram_do_i1_017 }),
    .f({\picorv32_core/cpuregs_rs2 [31],\picorv32_core/cpuregs_rs2 [17]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0100010001010000),
    .MODE("LOGIC"))
    \_al_u1363|_al_u1403  (
    .a({_al_u1308_o,_al_u1308_o}),
    .b({\picorv32_core/cpuregs_p2/dram_do_i1_030 ,\picorv32_core/decoded_rs2 [4]}),
    .c({\picorv32_core/cpuregs_p2/dram_do_i0_030 ,\picorv32_core/cpuregs_p2/dram_do_i0_018 }),
    .d({\picorv32_core/decoded_rs2 [4],\picorv32_core/cpuregs_p2/dram_do_i1_018 }),
    .f({\picorv32_core/cpuregs_rs2 [30],\picorv32_core/cpuregs_rs2 [18]}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~C*~B*~D+A*C*~B*~D+A*~C*B*~D+A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+A*C*B*D"),
    //.LUTF1("~B*A*~C*D+B*A*~C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG0("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG1("~B*A*C*~D+B*A*C*~D+~B*A*C*D+B*A*C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111110101010),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b1111111111111111),
    .INIT_LUTG1(16'b1010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1365|picorv32_core/reg26_b2  (
    .a({\picorv32_core/n664_lutinv_placeOpt_3 ,\picorv32_core/sel42_b2/B5 }),
    .c({\picorv32_core/cpuregs_rs2 [2],_al_u1339_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoded_imm [2],mem_la_wdata[2]}),
    .e({\picorv32_core/n523_lutinv ,\picorv32_core/sel42_b2/B4 }),
    .f({\picorv32_core/sel42_b2/B5 ,open_n5066}),
    .q({open_n5070,mem_la_wdata[2]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*~B)*~(D*C*~A))"),
    //.LUT1("(~(1*~B)*~(A*D*~C))"),
    .INIT_LUT0(16'b1010111111111111),
    .INIT_LUT1(16'b1100010011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1367 (
    .a({\picorv32_core/decoded_imm [29],\picorv32_core/n523_lutinv }),
    .b({_al_u1339_o,_al_u1339_o}),
    .c({\picorv32_core/n523_lutinv ,\picorv32_core/n664_lutinv_placeOpt_7 }),
    .d({\picorv32_core/n664_lutinv_placeOpt_7 ,\picorv32_core/decoded_imm [29]}),
    .mi({open_n5083,\picorv32_core/pcpi_rs2$29$ }),
    .fx({open_n5088,_al_u1367_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~A))"),
    //.LUT1("(~A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101111100001111),
    .INIT_LUT1(16'b0100010001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1368|picorv32_core/reg26_b29  (
    .a({_al_u1308_o,_al_u1337_o}),
    .b({\picorv32_core/cpuregs_p2/dram_do_i1_029 ,open_n5091}),
    .c({\picorv32_core/cpuregs_p2/dram_do_i0_029 ,_al_u1367_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoded_rs2 [4],\picorv32_core/cpuregs_rs2 [29]}),
    .f({\picorv32_core/cpuregs_rs2 [29],open_n5105}),
    .q({open_n5109,\picorv32_core/pcpi_rs2$29$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*~B)*~(D*C*~A))"),
    //.LUT1("(~(1*~B)*~(A*C*~D))"),
    .INIT_LUT0(16'b1010111111111111),
    .INIT_LUT1(16'b1100110001001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1370 (
    .a({\picorv32_core/decoded_imm [28],\picorv32_core/n523_lutinv }),
    .b({_al_u1339_o,_al_u1339_o}),
    .c({\picorv32_core/n664_lutinv_placeOpt_7 ,\picorv32_core/n664_lutinv_placeOpt_7 }),
    .d({\picorv32_core/n523_lutinv ,\picorv32_core/decoded_imm [28]}),
    .mi({open_n5122,\picorv32_core/pcpi_rs2$28$ }),
    .fx({open_n5127,_al_u1370_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~A))"),
    //.LUT1("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101111100001111),
    .INIT_LUT1(16'b0011001000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1371|picorv32_core/reg26_b28  (
    .a({\picorv32_core/cpuregs_p2/dram_do_i0_028 ,_al_u1337_o}),
    .b({_al_u1308_o,open_n5130}),
    .c({\picorv32_core/decoded_rs2 [4],_al_u1370_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_p2/dram_do_i1_028 ,\picorv32_core/cpuregs_rs2 [28]}),
    .f({\picorv32_core/cpuregs_rs2 [28],open_n5144}),
    .q({open_n5148,\picorv32_core/pcpi_rs2$28$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0011001000000010),
    .MODE("LOGIC"))
    \_al_u1374|_al_u1400  (
    .a({\picorv32_core/cpuregs_p2/dram_do_i0_027 ,_al_u1308_o}),
    .b({_al_u1308_o,\picorv32_core/decoded_rs2 [4]}),
    .c({\picorv32_core/decoded_rs2 [4],\picorv32_core/cpuregs_p2/dram_do_i0_019 }),
    .d({\picorv32_core/cpuregs_p2/dram_do_i1_027 ,\picorv32_core/cpuregs_p2/dram_do_i1_019 }),
    .f({\picorv32_core/cpuregs_rs2 [27],\picorv32_core/cpuregs_rs2 [19]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*C*~B*D+~A*C*B*D"),
    //.LUTF1("A*B*~C*~D+A*B*C*~D"),
    //.LUTG0("~A*~C*~B*~D+~A*~C*B*~D+~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    .INIT_LUTF0(16'b0101000000000000),
    .INIT_LUTF1(16'b0000000010001000),
    .INIT_LUTG0(16'b0101010100000101),
    .INIT_LUTG1(16'b0000000011011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1377|_al_u1392  (
    .a({\picorv32_core/decoded_rs2 [4],_al_u1308_o}),
    .b({\picorv32_core/cpuregs_p2/dram_do_i1_026 ,open_n5169}),
    .c({open_n5170,\picorv32_core/decoded_rs2 [4]}),
    .d({_al_u1308_o,\picorv32_core/cpuregs_p2/dram_do_i1_021 }),
    .e({\picorv32_core/cpuregs_p2/dram_do_i0_026 ,\picorv32_core/cpuregs_p2/dram_do_i0_021 }),
    .f({\picorv32_core/cpuregs_rs2 [26],\picorv32_core/cpuregs_rs2 [21]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*~B)*~(D*C*~A))"),
    //.LUT1("(~(1*~B)*~(A*C*~D))"),
    .INIT_LUT0(16'b1010111111111111),
    .INIT_LUT1(16'b1100110001001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1379 (
    .a({\picorv32_core/decoded_imm [25],\picorv32_core/n523_lutinv }),
    .b({_al_u1339_o,_al_u1339_o}),
    .c({\picorv32_core/n664_lutinv_placeOpt_6 ,\picorv32_core/n664_lutinv_placeOpt_6 }),
    .d({\picorv32_core/n523_lutinv ,\picorv32_core/decoded_imm [25]}),
    .mi({open_n5205,\picorv32_core/pcpi_rs2$25$ }),
    .fx({open_n5210,_al_u1379_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~A))"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*~C*D+A*B*~C*D"),
    //.LUTG0("~(C*~(D*~A))"),
    //.LUTG1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101111100001111),
    .INIT_LUTF1(16'b0000101000001010),
    .INIT_LUTG0(16'b0101111100001111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1380|picorv32_core/reg26_b25  (
    .a({\picorv32_core/cpuregs_p2/dram_do_i0_025 ,_al_u1337_o}),
    .c({_al_u1308_o,_al_u1379_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_p2/dram_do_i1_025 ,\picorv32_core/cpuregs_rs2 [25]}),
    .e({\picorv32_core/decoded_rs2 [4],open_n5215}),
    .f({\picorv32_core/cpuregs_rs2 [25],open_n5231}),
    .q({open_n5235,\picorv32_core/pcpi_rs2$25$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*~B)*~(D*C*~A))"),
    //.LUT1("(~(1*~B)*~(D*C*~A))"),
    .INIT_LUT0(16'b1010111111111111),
    .INIT_LUT1(16'b1000110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1382 (
    .a({\picorv32_core/n523_lutinv ,\picorv32_core/n523_lutinv }),
    .b({_al_u1339_o,_al_u1339_o}),
    .c({\picorv32_core/n664_lutinv_placeOpt_6 ,\picorv32_core/n664_lutinv_placeOpt_6 }),
    .d({\picorv32_core/decoded_imm [24],\picorv32_core/decoded_imm [24]}),
    .mi({open_n5248,\picorv32_core/pcpi_rs2$24$ }),
    .fx({open_n5253,_al_u1382_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D*~A))"),
    //.LUTF1("~B*A*~C*D+B*A*~C*D"),
    //.LUTG0("~(B*~(D*~A))"),
    //.LUTG1("~B*~A*~C*~D+B*~A*~C*~D+~B*~A*~C*D+B*~A*~C*D+~B*A*~C*D+B*A*~C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100110011),
    .INIT_LUTF1(16'b0000101000000000),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0000111100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1383|picorv32_core/reg26_b24  (
    .a({\picorv32_core/decoded_rs2 [4],_al_u1337_o}),
    .b({open_n5256,_al_u1382_o}),
    .c({_al_u1308_o,open_n5257}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_p2/dram_do_i1_024 ,\picorv32_core/cpuregs_rs2 [24]}),
    .e({\picorv32_core/cpuregs_p2/dram_do_i0_024 ,open_n5258}),
    .f({\picorv32_core/cpuregs_rs2 [24],open_n5274}),
    .q({open_n5278,\picorv32_core/pcpi_rs2$24$ }));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*B*~A*D+~C*B*A*D"),
    //.LUTF1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("~C*~B*~A*~D+~C*~B*A*~D+~C*~B*~A*D+~C*B*~A*D+~C*~B*A*D+~C*B*A*D"),
    //.LUTG1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000111000000010),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1386|_al_u1389  (
    .a({\picorv32_core/cpuregs_p2/dram_do_i0_023 ,open_n5279}),
    .b({\picorv32_core/decoded_rs2 [4],\picorv32_core/decoded_rs2 [4]}),
    .c({_al_u1308_o,_al_u1308_o}),
    .d({\picorv32_core/cpuregs_p2/dram_do_i1_023 ,\picorv32_core/cpuregs_p2/dram_do_i1_022 }),
    .e({open_n5282,\picorv32_core/cpuregs_p2/dram_do_i0_022 }),
    .f(\picorv32_core/cpuregs_rs2 [23:22]));
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*~B)*~(D*C*~A))"),
    //.LUT1("(~(1*~D)*~(B*C*~A))"),
    .INIT_LUT0(16'b1010111111111111),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1391 (
    .a({\picorv32_core/n523_lutinv ,\picorv32_core/n523_lutinv }),
    .b({\picorv32_core/decoded_imm [21],_al_u1339_o}),
    .c({\picorv32_core/n664_lutinv_placeOpt_1 ,\picorv32_core/n664_lutinv_placeOpt_1 }),
    .d({_al_u1339_o,\picorv32_core/decoded_imm [21]}),
    .mi({open_n5315,\picorv32_core/pcpi_rs2$21$ }),
    .fx({open_n5320,_al_u1391_o}));
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D"),
    //.LUTF1("(~(0*~C)*~(D*B*~A))"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("(~(1*~C)*~(D*B*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010101010),
    .INIT_LUTF1(16'b1011101111111111),
    .INIT_LUTG0(16'b1111111110101010),
    .INIT_LUTG1(16'b1011000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1394|uart/reg2_b20  (
    .a({\picorv32_core/n523_lutinv ,mem_la_wdata[4]}),
    .b({\picorv32_core/n664_lutinv_placeOpt_7 ,open_n5323}),
    .c({_al_u1339_o,open_n5324}),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\picorv32_core/decoded_imm [20],\picorv32_core/n734_lutinv }),
    .e({\picorv32_core/pcpi_rs2$20$ ,\picorv32_core/pcpi_rs2$20$ }),
    .sr(resetn_placeOpt_13),
    .f({_al_u1394_o,mem_la_wdata[20]}),
    .q({open_n5342,\uart/uart_bsrr [20]}));  // ../src/uart.v(102)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~A))"),
    //.LUT1("(~A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101111100001111),
    .INIT_LUT1(16'b0100010001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1395|picorv32_core/reg26_b20  (
    .a({_al_u1308_o,_al_u1337_o}),
    .b({\picorv32_core/cpuregs_p2/dram_do_i1_020 ,open_n5343}),
    .c({\picorv32_core/cpuregs_p2/dram_do_i0_020 ,_al_u1394_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoded_rs2 [4],\picorv32_core/cpuregs_rs2 [20]}),
    .f({\picorv32_core/cpuregs_rs2 [20],open_n5357}),
    .q({open_n5361,\picorv32_core/pcpi_rs2$20$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*~B)*~(D*C*~A))"),
    //.LUT1("(~(1*~D)*~(B*C*~A))"),
    .INIT_LUT0(16'b1010111111111111),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1399 (
    .a({\picorv32_core/n523_lutinv ,\picorv32_core/n523_lutinv }),
    .b({\picorv32_core/decoded_imm [19],_al_u1339_o}),
    .c({\picorv32_core/n664_lutinv_placeOpt_1 ,\picorv32_core/n664_lutinv_placeOpt_1 }),
    .d({_al_u1339_o,\picorv32_core/decoded_imm [19]}),
    .mi({open_n5374,\picorv32_core/pcpi_rs2$19$ }),
    .fx({open_n5379,_al_u1399_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*~B)*~(D*C*~A))"),
    //.LUT1("(~(1*~B)*~(D*C*~A))"),
    .INIT_LUT0(16'b1010111111111111),
    .INIT_LUT1(16'b1000110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1408 (
    .a({\picorv32_core/n523_lutinv ,\picorv32_core/n523_lutinv }),
    .b({_al_u1339_o,_al_u1339_o}),
    .c({\picorv32_core/n664_lutinv ,\picorv32_core/n664_lutinv }),
    .d({\picorv32_core/decoded_imm [16],\picorv32_core/decoded_imm [16]}),
    .mi({open_n5394,\picorv32_core/pcpi_rs2$16$ }),
    .fx({open_n5399,_al_u1408_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~A))"),
    //.LUT1("(~A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101111100001111),
    .INIT_LUT1(16'b0100010001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1409|picorv32_core/reg26_b16  (
    .a({_al_u1308_o,_al_u1337_o}),
    .b({\picorv32_core/cpuregs_p2/dram_do_i1_016 ,open_n5402}),
    .c({\picorv32_core/cpuregs_p2/dram_do_i0_016 ,_al_u1408_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoded_rs2 [4],\picorv32_core/cpuregs_rs2 [16]}),
    .f({\picorv32_core/cpuregs_rs2 [16],open_n5416}),
    .q({open_n5420,\picorv32_core/pcpi_rs2$16$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*~B)*~(D*C*~A))"),
    //.LUT1("(~(1*~B)*~(D*C*~A))"),
    .INIT_LUT0(16'b1010111111111111),
    .INIT_LUT1(16'b1000110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1414 (
    .a({\picorv32_core/n523_lutinv ,\picorv32_core/n523_lutinv }),
    .b({_al_u1339_o,_al_u1339_o}),
    .c({\picorv32_core/n664_lutinv ,\picorv32_core/n664_lutinv }),
    .d({\picorv32_core/decoded_imm [14],\picorv32_core/decoded_imm [14]}),
    .mi({open_n5433,\picorv32_core/pcpi_rs2$14$ }),
    .fx({open_n5438,_al_u1414_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D*~C))"),
    //.LUT1("(~A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100110011),
    .INIT_LUT1(16'b0100010001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1415|picorv32_core/reg26_b14  (
    .a({_al_u1308_o,open_n5441}),
    .b({\picorv32_core/cpuregs_p2/dram_do_i1_014 ,_al_u1414_o}),
    .c({\picorv32_core/cpuregs_p2/dram_do_i0_014 ,_al_u1337_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoded_rs2 [4],\picorv32_core/cpuregs_rs2 [14]}),
    .f({\picorv32_core/cpuregs_rs2 [14],open_n5455}),
    .q({open_n5459,\picorv32_core/pcpi_rs2$14$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*~B)*~(D*C*~A))"),
    //.LUT1("(~(1*~B)*~(A*D*~C))"),
    .INIT_LUT0(16'b1010111111111111),
    .INIT_LUT1(16'b1100010011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1417 (
    .a({\picorv32_core/decoded_imm [13],\picorv32_core/n523_lutinv }),
    .b({_al_u1339_o,_al_u1339_o}),
    .c({\picorv32_core/n523_lutinv ,\picorv32_core/n664_lutinv }),
    .d({\picorv32_core/n664_lutinv ,\picorv32_core/decoded_imm [13]}),
    .mi({open_n5472,\picorv32_core/pcpi_rs2$13$ }),
    .fx({open_n5477,_al_u1417_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~(D*~C))"),
    //.LUTF1("A*~B*~D*~C+A*~B*~D*C"),
    //.LUTG0("~(A*~(D*~C))"),
    //.LUTG1("A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101111101010101),
    .INIT_LUTF1(16'b0000000000100010),
    .INIT_LUTG0(16'b0101111101010101),
    .INIT_LUTG1(16'b0000000011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1418|picorv32_core/reg26_b13  (
    .a({\picorv32_core/cpuregs_p2/dram_do_i0_013 ,_al_u1417_o}),
    .b({\picorv32_core/decoded_rs2 [4],open_n5480}),
    .c({open_n5481,_al_u1337_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1308_o,\picorv32_core/cpuregs_rs2 [13]}),
    .e({\picorv32_core/cpuregs_p2/dram_do_i1_013 ,open_n5482}),
    .f({\picorv32_core/cpuregs_rs2 [13],open_n5498}),
    .q({open_n5502,\picorv32_core/pcpi_rs2$13$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*~B)*~(D*C*~A))"),
    //.LUT1("(~(1*~D)*~(B*C*~A))"),
    .INIT_LUT0(16'b1010111111111111),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1426 (
    .a({\picorv32_core/n523_lutinv ,\picorv32_core/n523_lutinv }),
    .b({\picorv32_core/decoded_imm [10],_al_u1339_o}),
    .c({\picorv32_core/n664_lutinv_placeOpt_7 ,\picorv32_core/n664_lutinv_placeOpt_7 }),
    .d({_al_u1339_o,\picorv32_core/decoded_imm [10]}),
    .mi({open_n5515,\picorv32_core/pcpi_rs2$10$ }),
    .fx({open_n5520,_al_u1426_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D*~A))"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*~C*D+A*B*~C*D"),
    //.LUTG0("~(B*~(D*~A))"),
    //.LUTG1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100110011),
    .INIT_LUTF1(16'b0000101000001010),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1427|picorv32_core/reg26_b10  (
    .a({\picorv32_core/cpuregs_p2/dram_do_i0_010 ,_al_u1337_o}),
    .b({open_n5523,_al_u1426_o}),
    .c({_al_u1308_o,open_n5524}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_p2/dram_do_i1_010 ,\picorv32_core/cpuregs_rs2 [10]}),
    .e({\picorv32_core/decoded_rs2 [4],open_n5525}),
    .f({\picorv32_core/cpuregs_rs2 [10],open_n5541}),
    .q({open_n5545,\picorv32_core/pcpi_rs2$10$ }));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101110101010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111111111111111),
    .INIT_LUTG1(16'b1101100011011000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1429|picorv32_core/reg26_b0  (
    .a({\picorv32_core/n523_lutinv ,\picorv32_core/sel42_b0/B5 }),
    .b({\picorv32_core/cpuregs_rs2 [0],_al_u1339_o}),
    .c({\picorv32_core/decoded_imm [0],open_n5546}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({open_n5547,mem_la_wdata[0]}),
    .e({\picorv32_core/n664_lutinv_placeOpt_6 ,\picorv32_core/sel42_b0/B4 }),
    .f({\picorv32_core/sel42_b0/B5 ,open_n5563}),
    .q({open_n5567,mem_la_wdata[0]}));  // ../src/picorv32.v(1906)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~D*~C*~B*~A+D*~C*~B*~A+~D*C*~B*~A+D*C*~B*~A+~D*~C*B*~A+D*~C*B*~A+~D*C*B*~A+~D*C*~B*A+D*C*~B*A+~D*C*B*A"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~D*~C*~B*~A+D*~C*~B*~A+D*C*~B*~A+~D*~C*B*~A+D*~C*B*~A+D*C*~B*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0011010111110101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0011010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1431|uart/reg0_b14  (
    .a({\picorv32_core/mem_rdata_q [14],\picorv32_core/pcpi_rs1$3$ }),
    .b({uart_do[14],\picorv32_core/n30 [1]}),
    .c({\picorv32_core/mem_xfer_placeOpt_4 ,_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_2,mem_la_addr[2]}),
    .e({memory_out[14],\uart/uart_bsrr [14]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1431_o,open_n5582}),
    .q({open_n5586,uart_do[14]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("~D*~C*~B*~A+D*~C*~B*~A+~D*C*~B*~A+D*C*~B*~A+~D*~C*B*~A+D*~C*B*~A+~D*C*B*~A+D*C*B*~A"),
    //.LUTG0("(1*~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("~D*~C*~B*~A+D*~C*~B*~A+D*C*~B*~A+~D*~C*B*~A+~D*~C*~B*A+D*~C*~B*A+D*C*~B*A+~D*~C*B*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000000011001010),
    .INIT_LUTG1(16'b0011001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1432|uart/reg0_b30  (
    .a({\picorv32_core/mem_rdata_q [30],\picorv32_core/n30 [1]}),
    .b({uart_do[30],\picorv32_core/pcpi_rs1$3$ }),
    .c({memory_out[30],_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_2,mem_la_addr[2]}),
    .e({\picorv32_core/mem_xfer_placeOpt_4 ,\uart/uart_bsrr [30]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1432_o,open_n5601}),
    .q({open_n5605,uart_do[30]}));  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*~B)"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"))
    \_al_u1433|_al_u1258  (
    .a({\picorv32_core/mem_la_secondword ,\picorv32_core/mem_la_secondword }),
    .b({_al_u1088_o,open_n5606}),
    .d({open_n5611,_al_u1089_o}),
    .f({\picorv32_core/mux3_b16_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG0("~(~1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+~A*~B*C*D"),
    .INIT_LUTF0(16'b0000001010001010),
    .INIT_LUTF1(16'b0001000100000011),
    .INIT_LUTG0(16'b0101011111011111),
    .INIT_LUTG1(16'b0001000100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1434|_al_u1483  (
    .a({_al_u1432_o,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({_al_u1089_o,_al_u1088_o}),
    .c({_al_u1431_o,_al_u1431_o}),
    .d({\picorv32_core/mux3_b16_sel_is_0_o ,_al_u1432_o}),
    .e({open_n5632,\picorv32_core/mem_16bit_buffer [14]}),
    .f({\picorv32_core/mem_rdata_latched [30],_al_u1483_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*~B*~D*~C+A*~B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*~B*~D*C+~A*B*~D*C+~A*~B*D*C+~A*B*D*C"),
    //.LUTG0("~(~1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000001010001010),
    .INIT_LUTF1(16'b0101001101010011),
    .INIT_LUTG0(16'b0101011111011111),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1434|_al_u1483_placeOpt_1  (
    .a({_al_u1432_o,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({_al_u1431_o,_al_u1088_o}),
    .c({\picorv32_core/mux3_b16_sel_is_0_o ,_al_u1431_o}),
    .d({open_n5655,_al_u1432_o}),
    .e({_al_u1089_o,\picorv32_core/mem_16bit_buffer [14]}),
    .f({open_n5671,_al_u1483_o_placeOpt_1}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*~B*D+~A*C*~B*D"),
    //.LUTG0("~(~1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*~C*~B*D+~A*C*~B*D"),
    .INIT_LUTF0(16'b0000001010001010),
    .INIT_LUTF1(16'b0001000100110011),
    .INIT_LUTG0(16'b0101011111011111),
    .INIT_LUTG1(16'b0001000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1434|_al_u1483_placeOpt_2  (
    .a({_al_u1432_o,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({_al_u1089_o,_al_u1088_o}),
    .c({open_n5677,_al_u1431_o}),
    .d({\picorv32_core/mux3_b16_sel_is_0_o ,_al_u1432_o}),
    .e({_al_u1431_o,\picorv32_core/mem_16bit_buffer [14]}),
    .f({open_n5695,_al_u1483_o_placeOpt_2}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~(~1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000001010001010),
    .INIT_LUTF1(16'b0101010100110011),
    .INIT_LUTG0(16'b0101011111011111),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1434|_al_u1483_placeOpt_3  (
    .a({_al_u1432_o,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({_al_u1431_o,_al_u1088_o}),
    .c({open_n5701,_al_u1431_o}),
    .d({\picorv32_core/mux3_b16_sel_is_0_o ,_al_u1432_o}),
    .e({_al_u1089_o,\picorv32_core/mem_16bit_buffer [14]}),
    .f({open_n5719,_al_u1483_o_placeOpt_3}));
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~(A*~((B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D))*~(C)+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*~(C)+~(A)*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C)"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~(A*~((B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D))*~(C)+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*~(C)+~(A)*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111010100110101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0000010100110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1435|uart/reg0_b24  (
    .a({\picorv32_core/mem_rdata_q [24],\picorv32_core/pcpi_rs1$3$ }),
    .b({memory_out[24],\picorv32_core/n30 [1]}),
    .c({\picorv32_core/mem_xfer_placeOpt_5 ,_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_3,mem_la_addr[2]}),
    .e({uart_do[24],\uart/uart_bsrr [24]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1435_o,open_n5739}),
    .q({open_n5743,uart_do[24]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~(B*~((A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C))*~(D)+B*(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*~(D)+~(B)*(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*D+B*(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*D)"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~(B*~((A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C))*~(D)+B*(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*~(D)+~(B)*(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*D+B*(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111010100110011),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0000010100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1436|uart/reg0_b8  (
    .a({memory_out[8],\picorv32_core/pcpi_rs1$3$ }),
    .b({\picorv32_core/mem_rdata_q [8],\picorv32_core/n30 [1]}),
    .c({uart_sel_lutinv_placeOpt_3,_al_u700_o_placeOpt_2}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_xfer_placeOpt_5 ,mem_la_addr[2]}),
    .e({uart_do[8],\uart/uart_bsrr [8]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1436_o,open_n5758}),
    .q({open_n5762,uart_do[8]}));  // ../src/uart.v(102)
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~D*~C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+A*~D*~C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    //.LUTF1("A*~D*~C*~B+A*~D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+~A*~D*C*B+A*~D*C*B+~A*D*C*B"),
    //.LUTG0("~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+A*~D*~C*B+A*D*~C*B+A*~D*C*B+A*D*C*B"),
    //.LUTG1("A*~D*~C*~B+A*D*~C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+~A*D*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000010101010),
    .INIT_LUTF1(16'b0100010011101110),
    .INIT_LUTG0(16'b1011100010111000),
    .INIT_LUTG1(16'b0100111001001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1437|picorv32_core/reg5_b8  (
    .a({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mem_16bit_buffer [8]}),
    .b({\picorv32_core/mem_16bit_buffer [8],_al_u1089_o}),
    .c({_al_u1435_o,mem_rdata[24]}),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u1436_o,\picorv32_core/mux51_b0_sel_is_3_o }),
    .e({_al_u1088_o,\picorv32_core/mem_la_read }),
    .f({\picorv32_core/mux79_b1/B0_3 ,open_n5778}),
    .q({open_n5782,\picorv32_core/mem_16bit_buffer [8]}));  // ../src/picorv32.v(605)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~(A*~((B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D))*~(C)+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*~(C)+~(A)*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C)"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~(A*~((B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D))*~(C)+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*~(C)+~(A)*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111010100110101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0000010100110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1439|uart/reg0_b13  (
    .a({\picorv32_core/mem_rdata_q [13],\picorv32_core/pcpi_rs1$3$ }),
    .b({memory_out[13],\picorv32_core/n30 [1]}),
    .c({\picorv32_core/mem_xfer ,_al_u700_o_placeOpt_2}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_3,mem_la_addr[2]}),
    .e({uart_do[13],\uart/uart_bsrr [13]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1439_o,open_n5797}),
    .q({open_n5801,uart_do[13]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*~B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0011001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1440|uart/reg0_b29  (
    .a({\picorv32_core/mem_rdata_q [29],\picorv32_core/pcpi_rs1$3$ }),
    .b({uart_do[29],\picorv32_core/n30 [1]}),
    .c({memory_out[29],_al_u700_o_placeOpt_2}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_2,mem_la_addr[2]}),
    .e({\picorv32_core/mem_xfer ,\uart/uart_bsrr [29]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1440_o,open_n5816}),
    .q({open_n5820,uart_do[29]}));  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*D*~C+B*~A*D*~C+~B*A*D*~C+B*A*D*~C+~B*~A*D*C+B*~A*D*C+~B*A*D*C+B*A*D*C"),
    //.LUTF1("~A*~C*~D*~B+A*~C*~D*~B+~A*C*~D*~B+A*C*~D*~B+~A*C*D*~B+A*C*D*~B+~A*~C*~D*B+A*~C*~D*B"),
    //.LUTG0("~B*~A*D*C+B*~A*D*C+~B*A*D*C+B*A*D*C"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1441|_al_u1637  (
    .b({_al_u1440_o,open_n5823}),
    .c({\picorv32_core/mux3_b16_sel_is_0_o ,_al_u1440_o}),
    .d({_al_u1439_o,\picorv32_core/mux4_b0_sel_is_0_o }),
    .e({_al_u1089_o,_al_u1088_o}),
    .f({\picorv32_core/mem_rdata_latched [29],_al_u1637_o}));
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*~B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0011001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1442|uart/reg0_b10  (
    .a({\picorv32_core/mem_rdata_q [10],\picorv32_core/pcpi_rs1$3$ }),
    .b({uart_do[10],\picorv32_core/n30 [1]}),
    .c({memory_out[10],_al_u700_o_placeOpt_2}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_3,mem_la_addr[2]}),
    .e({\picorv32_core/mem_xfer_placeOpt_5 ,\uart/uart_bsrr [10]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1442_o,open_n5860}),
    .q({open_n5864,uart_do[10]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~(B*~((A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C))*~(D)+B*(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*~(D)+~(B)*(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*D+B*(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*D)"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~(B*~((A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C))*~(D)+B*(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*~(D)+~(B)*(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*D+B*(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111010100110011),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0000010100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1443|uart/reg0_b26  (
    .a({memory_out[26],\picorv32_core/pcpi_rs1$3$ }),
    .b({\picorv32_core/mem_rdata_q [26],\picorv32_core/n30 [1]}),
    .c({uart_sel_lutinv_placeOpt_3,_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_xfer_placeOpt_5 ,mem_la_addr[2]}),
    .e({uart_do[26],\uart/uart_bsrr [26]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1443_o,open_n5879}),
    .q({open_n5883,uart_do[26]}));  // ../src/uart.v(102)
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~D*~C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+A*~D*~C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    //.LUTF1("~D*~C*B*~A+~D*C*B*~A+~D*~C*~B*A+D*~C*~B*A+~D*C*~B*A+D*C*~B*A+~D*~C*B*A+~D*C*B*A"),
    //.LUTG0("~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+A*~D*~C*B+A*D*~C*B+A*~D*C*B+A*D*C*B"),
    //.LUTG1("~D*~C*B*~A+D*~C*B*~A+~D*~C*~B*A+D*~C*~B*A+~D*C*~B*A+D*C*~B*A+~D*~C*B*A+D*~C*B*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000010101010),
    .INIT_LUTF1(16'b0010001011101110),
    .INIT_LUTG0(16'b1011100010111000),
    .INIT_LUTG1(16'b0010111000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1444|picorv32_core/reg5_b10  (
    .a({\picorv32_core/mem_16bit_buffer [10],\picorv32_core/mem_16bit_buffer [10]}),
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,_al_u1089_o}),
    .c({_al_u1443_o,mem_rdata[26]}),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u1442_o,\picorv32_core/mux51_b0_sel_is_3_o }),
    .e({_al_u1088_o,\picorv32_core/mem_la_read }),
    .f({_al_u1444_o,open_n5899}),
    .q({open_n5903,\picorv32_core/mem_16bit_buffer [10]}));  // ../src/picorv32.v(605)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~0*~((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))*~(A)+~0*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*~(A)+~(~0)*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*A+~0*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*A)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*~C*D+A*B*~C*D"),
    //.LUTG0("~(~1*~((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))*~(A)+~1*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*~(A)+~(~1)*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*A+~1*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*A)"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000101010),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0101110101111111),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1446|picorv32_core/reg6_b12  (
    .a({open_n5904,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({\picorv32_core/mux3_b16_sel_is_0_o ,_al_u1088_o}),
    .c({_al_u1272_o,_al_u1272_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u1273_o,_al_u1273_o}),
    .e({_al_u1089_o,\picorv32_core/mem_16bit_buffer [12]}),
    .f({\picorv32_core/mem_rdata_latched [28],\picorv32_core/mem_rdata_latched [12]}),
    .q({open_n5923,\picorv32_core/decoded_imm_uj [12]}));  // ../src/picorv32.v(1120)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    //.LUTG0("(1*~A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*~B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0101010000000100),
    .INIT_LUTG1(16'b0011001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1447|uart/reg0_b9  (
    .a({\picorv32_core/mem_rdata_q [9],mem_la_addr[2]}),
    .b({uart_do[9],\picorv32_core/n30 [1]}),
    .c({memory_out[9],_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_3,\picorv32_core/pcpi_rs1$3$ }),
    .e({\picorv32_core/mem_xfer_placeOpt_5 ,\uart/uart_bsrr [9]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1447_o,open_n5938}),
    .q({open_n5942,uart_do[9]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~(B*~((A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C))*~(D)+B*(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*~(D)+~(B)*(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*D+B*(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*D)"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~(B*~((A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C))*~(D)+B*(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*~(D)+~(B)*(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*D+B*(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111010100110011),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0000010100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1448|uart/reg0_b25  (
    .a({memory_out[25],\picorv32_core/pcpi_rs1$3$ }),
    .b({\picorv32_core/mem_rdata_q [25],\picorv32_core/n30 [1]}),
    .c({uart_sel_lutinv_placeOpt_2,_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_xfer_placeOpt_4 ,mem_la_addr[2]}),
    .e({uart_do[25],\uart/uart_bsrr [25]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1448_o,open_n5957}),
    .q({open_n5961,uart_do[25]}));  // ../src/uart.v(102)
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~D*~C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+A*~D*~C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    //.LUTF1("~D*B*~C*~A+~D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A"),
    //.LUTG0("~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+A*~D*~C*B+A*D*~C*B+A*~D*C*B+A*D*C*B"),
    //.LUTG1("~D*B*~C*~A+D*B*~C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+D*~B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000010101010),
    .INIT_LUTF1(16'b0010001011101110),
    .INIT_LUTG0(16'b1011100010111000),
    .INIT_LUTG1(16'b0010111000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1449|picorv32_core/reg5_b9  (
    .a({\picorv32_core/mem_16bit_buffer [9],\picorv32_core/mem_16bit_buffer [9]}),
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,_al_u1089_o}),
    .c({_al_u1448_o,mem_rdata[25]}),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u1447_o,\picorv32_core/mux51_b0_sel_is_3_o }),
    .e({_al_u1088_o,\picorv32_core/mem_la_read }),
    .f({\picorv32_core/mux79_b2/B0_3 ,open_n5977}),
    .q({open_n5981,\picorv32_core/mem_16bit_buffer [9]}));  // ../src/picorv32.v(605)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*~B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0011001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1451|uart/reg0_b11  (
    .a({\picorv32_core/mem_rdata_q [11],\picorv32_core/pcpi_rs1$3$ }),
    .b({uart_do[11],\picorv32_core/n30 [1]}),
    .c({memory_out[11],_al_u700_o_placeOpt_2}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_3,mem_la_addr[2]}),
    .e({\picorv32_core/mem_xfer_placeOpt_5 ,\uart/uart_bsrr [11]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1451_o,open_n5996}),
    .q({open_n6000,uart_do[11]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~(A*~((B*~(0)*~(C)+B*0*~(C)+~(B)*0*C+B*0*C))*~(D)+A*(B*~(0)*~(C)+B*0*~(C)+~(B)*0*C+B*0*C)*~(D)+~(A)*(B*~(0)*~(C)+B*0*~(C)+~(B)*0*C+B*0*C)*D+A*(B*~(0)*~(C)+B*0*~(C)+~(B)*0*C+B*0*C)*D)"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~(A*~((B*~(1)*~(C)+B*1*~(C)+~(B)*1*C+B*1*C))*~(D)+A*(B*~(1)*~(C)+B*1*~(C)+~(B)*1*C+B*1*C)*~(D)+~(A)*(B*~(1)*~(C)+B*1*~(C)+~(B)*1*C+B*1*C)*D+A*(B*~(1)*~(C)+B*1*~(C)+~(B)*1*C+B*1*C)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111001101010101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0000001101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1452|uart/reg0_b27  (
    .a({\picorv32_core/mem_rdata_q [27],\picorv32_core/pcpi_rs1$3$ }),
    .b({memory_out[27],\picorv32_core/n30 [1]}),
    .c({uart_sel_lutinv_placeOpt_3,_al_u700_o_placeOpt_2}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_xfer_placeOpt_5 ,mem_la_addr[2]}),
    .e({uart_do[27],\uart/uart_bsrr [27]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1452_o,open_n6015}),
    .q({open_n6019,uart_do[27]}));  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D"),
    //.LUTG0("~(~1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000001010001010),
    .INIT_LUTF1(16'b0000001111001111),
    .INIT_LUTG0(16'b0101011111011111),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1453|_al_u1464  (
    .a({open_n6020,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({\picorv32_core/mux3_b16_sel_is_0_o ,_al_u1088_o}),
    .c({_al_u1451_o,_al_u1451_o}),
    .d({_al_u1452_o,_al_u1452_o}),
    .e({_al_u1089_o,\picorv32_core/mem_16bit_buffer [11]}),
    .f({\picorv32_core/mem_rdata_latched [27],_al_u1464_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0)*~((A*D*C))+B*0*~((A*D*C))+~(B)*0*(A*D*C)+B*0*(A*D*C))"),
    //.LUT1("(B*~(1)*~((A*D*C))+B*1*~((A*D*C))+~(B)*1*(A*D*C)+B*1*(A*D*C))"),
    .INIT_LUT0(16'b0100110011001100),
    .INIT_LUT1(16'b1110110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1455 (
    .a({_al_u1175_o,_al_u1175_o}),
    .b({memory_out[26],memory_out[26]}),
    .c({_al_u1279_o,_al_u1279_o}),
    .d({_al_u1168_o,_al_u1168_o}),
    .mi({open_n6055,uart_do[26]}),
    .fx({open_n6060,mem_rdata[26]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(0*~(D)*~(B)+0*D*~(B)+~(0)*D*B+0*D*B)))"),
    //.LUT1("(~A*~(D*~(1*~(C)*~(B)+1*C*~(B)+~(1)*C*B+1*C*B)))"),
    .INIT_LUT0(16'b0100010100000101),
    .INIT_LUT1(16'b0101000101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1456 (
    .a({_al_u1089_o,_al_u1089_o}),
    .b({\picorv32_core/mem_xfer_placeOpt_5 ,\picorv32_core/mem_xfer_placeOpt_5 }),
    .c({mem_rdata[26],\picorv32_core/mux3_b16_sel_is_0_o }),
    .d({\picorv32_core/mux3_b16_sel_is_0_o ,mem_rdata[26]}),
    .mi({open_n6075,\picorv32_core/mem_rdata_q [26]}),
    .fx({open_n6080,_al_u1456_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((D*~(~B*A)))*~(C)+0*(D*~(~B*A))*~(C)+~(0)*(D*~(~B*A))*C+0*(D*~(~B*A))*C)"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(1*~((D*~(~B*A)))*~(C)+1*(D*~(~B*A))*~(C)+~(1)*(D*~(~B*A))*C+1*(D*~(~B*A))*C)"),
    //.LUTG1("(B*~(~C*D))"),
    .INIT_LUTF0(16'b1101000000000000),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b1101111100001111),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1457|_al_u2409  (
    .a({open_n6083,_al_u1442_o}),
    .b({_al_u1456_o,\picorv32_core/mux3_b16_sel_is_0_o }),
    .c({\picorv32_core/mux3_b16_sel_is_0_o ,\picorv32_core/mem_xfer }),
    .d({_al_u1442_o,_al_u1456_o}),
    .e({open_n6086,\picorv32_core/mem_rdata_q [26]}),
    .f({\picorv32_core/mem_rdata_latched [26],\picorv32_core/n42 [26]}));
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*B*~(A)*~(0)+~(D)*~(C)*~(B)*A*~(0)+~(D)*~(C)*B*A*~(0)+D*~(C)*B*A*~(0)+~(D)*C*~(B)*~(A)*0+D*~(C)*B*~(A)*0+~(D)*C*B*~(A)*0+~(D)*~(C)*~(B)*A*0+~(D)*C*~(B)*A*0+~(D)*~(C)*B*A*0+D*~(C)*B*A*0+~(D)*C*B*A*0)"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    //.LUTG0("(D*~(C)*B*~(A)*~(1)+~(D)*~(C)*~(B)*A*~(1)+~(D)*~(C)*B*A*~(1)+D*~(C)*B*A*~(1)+~(D)*C*~(B)*~(A)*1+D*~(C)*B*~(A)*1+~(D)*C*B*~(A)*1+~(D)*~(C)*~(B)*A*1+~(D)*C*~(B)*A*1+~(D)*~(C)*B*A*1+D*~(C)*B*A*1+~(D)*C*B*A*1)"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*~B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110000001010),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000110011111010),
    .INIT_LUTG1(16'b0011001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1458|uart/reg0_b7  (
    .a({\picorv32_core/mem_rdata_q [7],\uart/uart_odr [7]}),
    .b({uart_do[7],\uart/uart_bsrr [7]}),
    .c({memory_out[7],mem_la_addr[2]}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_3,mem_la_addr[3]}),
    .e({\picorv32_core/mem_xfer_placeOpt_5 ,\uart/uart_idr [7]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1458_o,open_n6121}),
    .q({open_n6125,uart_do[7]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~(A*~((B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D))*~(C)+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*~(C)+~(A)*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C)"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~(A*~((B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D))*~(C)+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*~(C)+~(A)*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111010100110101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0000010100110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1459|uart/reg0_b23  (
    .a({\picorv32_core/mem_rdata_q [23],\picorv32_core/pcpi_rs1$3$ }),
    .b({memory_out[23],\picorv32_core/n30 [1]}),
    .c({\picorv32_core/mem_xfer_placeOpt_4 ,_al_u700_o_placeOpt_2}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_2,mem_la_addr[2]}),
    .e({uart_do[23],\uart/uart_bsrr [23]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1459_o,open_n6140}),
    .q({open_n6144,uart_do[23]}));  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUT1("~(~1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    .INIT_LUT0(16'b0000001010001010),
    .INIT_LUT1(16'b0101011111011111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1460 (
    .a({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({_al_u1088_o,_al_u1088_o}),
    .c({_al_u1458_o,_al_u1458_o}),
    .d({_al_u1459_o,_al_u1459_o}),
    .mi({open_n6157,\picorv32_core/mem_16bit_buffer [7]}),
    .fx({open_n6162,\picorv32_core/mux79_b0/B0_3 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*B)"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT_LUT0(16'b0100010001000100),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"))
    \_al_u1462|_al_u1500  (
    .a({\picorv32_core/mux3_b16_sel_is_0_o ,\picorv32_core/mem_do_rdata }),
    .b({_al_u1089_o,\picorv32_core/n131 }),
    .c({_al_u1448_o,open_n6165}),
    .d({_al_u1447_o,open_n6168}),
    .f({\picorv32_core/mem_rdata_latched [25],\picorv32_core/mux51_b0_sel_is_3_o }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUT0(16'b0000011100000100),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"))
    \_al_u1465|_al_u1491  (
    .a({_al_u1089_o,_al_u1261_o}),
    .b({\picorv32_core/mux3_b16_sel_is_0_o ,\picorv32_core/mux3_b16_sel_is_0_o }),
    .c({_al_u1436_o,_al_u1089_o}),
    .d({_al_u1435_o,\picorv32_core/mem_rdata_latched_noshuffle [5]}),
    .f({\picorv32_core/mem_rdata_latched [24],\picorv32_core/mem_rdata_latched [21]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUT0(16'b0000001111110011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"))
    \_al_u1467|_al_u2327  (
    .a({\picorv32_core/mux3_b16_sel_is_0_o ,open_n6207}),
    .b({_al_u1089_o,\picorv32_core/mem_rdata_q [23]}),
    .c({_al_u1458_o,\picorv32_core/mem_xfer }),
    .d({_al_u1459_o,\picorv32_core/mem_rdata_latched [23]}),
    .f({\picorv32_core/mem_rdata_latched [23],_al_u2327_o}));
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~(A*~((B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D))*~(C)+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*~(C)+~(A)*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C)"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~(A*~((B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D))*~(C)+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*~(C)+~(A)*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111010100110101),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0000010100110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1469|uart/reg0_b15  (
    .a({\picorv32_core/mem_rdata_q [15],\picorv32_core/pcpi_rs1$3$ }),
    .b({memory_out[15],\picorv32_core/n30 [1]}),
    .c({\picorv32_core/mem_xfer_placeOpt_4 ,_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_2,mem_la_addr[2]}),
    .e({uart_do[15],\uart/uart_bsrr [15]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1469_o,open_n6242}),
    .q({open_n6246,uart_do[15]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+~A*~D*C*B+A*~D*C*B"),
    //.LUTG0("(1*~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~A*D*~C*~B+~A*D*C*~B+A*D*C*~B+~A*D*~C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0011010111111111),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0011010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1470|uart/reg0_b31  (
    .a({memory_out[31],\picorv32_core/pcpi_rs1$3$ }),
    .b({uart_do[31],\picorv32_core/n30 [1]}),
    .c({uart_sel_lutinv_placeOpt_2,_al_u700_o_placeOpt_3}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_xfer_placeOpt_4 ,mem_la_addr[2]}),
    .e({\picorv32_core/mem_rdata_q [31],\uart/uart_bsrr [31]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1470_o,open_n6261}),
    .q({open_n6265,uart_do[31]}));  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT_LUT0(16'b0001001100000010),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"))
    \_al_u1471|_al_u1477  (
    .a({\picorv32_core/mux3_b16_sel_is_0_o ,\picorv32_core/mux3_b16_sel_is_0_o }),
    .b({_al_u1089_o,_al_u1089_o}),
    .c({_al_u1470_o,_al_u1276_o}),
    .d({_al_u1469_o,\picorv32_core/mem_rdata_latched_noshuffle [1]}),
    .f({\picorv32_core/mem_rdata_latched [31],\picorv32_core/mem_rdata_latched [17]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))"),
    //.LUT1("(~B*~(~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A))"),
    .INIT_LUT0(16'b0001001100000010),
    .INIT_LUT1(16'b0001000000110010),
    .MODE("LOGIC"))
    \_al_u1473|_al_u1489  (
    .a({\picorv32_core/mux3_b16_sel_is_0_o ,\picorv32_core/mux3_b16_sel_is_0_o }),
    .b({_al_u1089_o,_al_u1089_o}),
    .c({\picorv32_core/mem_rdata_latched_noshuffle [3],_al_u1257_o}),
    .d({_al_u1266_o,\picorv32_core/mem_rdata_latched_noshuffle [6]}),
    .f({\picorv32_core/mem_rdata_latched [19],\picorv32_core/mem_rdata_latched [22]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~B*D*~C*~A+B*D*~C*~A+~B*~D*C*~A+B*~D*C*~A+~B*D*C*~A+B*D*C*~A+~B*~D*C*A+B*~D*C*A"),
    //.LUTG0("~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0101010101000100),
    .INIT_LUTF1(16'b0101010111110000),
    .INIT_LUTG0(16'b0001000100000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1475|_al_u1487  (
    .a({_al_u1270_o,_al_u1089_o}),
    .b({open_n6306,\picorv32_core/mux3_b16_sel_is_0_o }),
    .c({\picorv32_core/mem_rdata_latched_noshuffle [2],open_n6307}),
    .d({\picorv32_core/mux3_b16_sel_is_0_o ,\picorv32_core/mem_rdata_latched_noshuffle [4]}),
    .e({_al_u1089_o,_al_u1264_o}),
    .f({\picorv32_core/mem_rdata_latched [18],\picorv32_core/mem_rdata_latched [20]}));
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTF1("~(~0*~((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))*~(A)+~0*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*~(A)+~(~0)*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*A+~0*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*A)"),
    //.LUTG0("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTG1("~(~1*~((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))*~(A)+~1*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*~(A)+~(~1)*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*A+~1*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010011000000),
    .INIT_LUTF1(16'b0000100000101010),
    .INIT_LUTG0(16'b1110111011001111),
    .INIT_LUTG1(16'b0101110101111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1481|picorv32_core/reg5_b15  (
    .a({\picorv32_core/mux4_b0_sel_is_0_o ,_al_u1089_o}),
    .b({_al_u1088_o,mem_rdata[31]}),
    .c({_al_u1470_o,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u1469_o,\picorv32_core/mem_la_read }),
    .e({\picorv32_core/mem_16bit_buffer [15],\picorv32_core/mem_16bit_buffer [15]}),
    .f({_al_u1481_o,open_n6345}),
    .q({open_n6349,\picorv32_core/mem_16bit_buffer [15]}));  // ../src/picorv32.v(605)
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTF1("~(~0*~((D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))*~(B)+~0*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*~(B)+~(~0)*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*B+~0*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*B)"),
    //.LUTG0("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTG1("~(~1*~((D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))*~(B)+~1*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*~(B)+~(~1)*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*B+~1*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010011000000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1110111011001111),
    .INIT_LUTG1(16'b0011101101111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1481|picorv32_core/reg5_b15_placeOpt_1  (
    .a({_al_u1088_o,_al_u1089_o}),
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,mem_rdata[31]}),
    .c({_al_u1470_o,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u1469_o,\picorv32_core/mem_la_read }),
    .e({\picorv32_core/mem_16bit_buffer [15],\picorv32_core/mem_16bit_buffer [15]}),
    .f({_al_u1481_o_placeOpt_1,open_n6365}));  // ../src/picorv32.v(605)
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTF1("~(~0*~((A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))*~(C)+~0*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)*~(C)+~(~0)*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)*C+~0*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)*C)"),
    //.LUTG0("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTG1("~(~1*~((A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))*~(C)+~1*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)*~(C)+~(~1)*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)*C+~1*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010011000000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1110111011001111),
    .INIT_LUTG1(16'b0001111111011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1481|picorv32_core/reg5_b15_placeOpt_2  (
    .a({_al_u1469_o,_al_u1089_o}),
    .b({_al_u1088_o,mem_rdata[31]}),
    .c({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u1470_o,\picorv32_core/mem_la_read }),
    .e({\picorv32_core/mem_16bit_buffer [15],\picorv32_core/mem_16bit_buffer [15]}),
    .f({_al_u1481_o_placeOpt_2,open_n6386}));  // ../src/picorv32.v(605)
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTF1("~(~0*~((D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))*~(B)+~0*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*~(B)+~(~0)*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*B+~0*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*B)"),
    //.LUTG0("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTG1("~(~1*~((D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))*~(B)+~1*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*~(B)+~(~1)*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*B+~1*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010011000000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1110111011001111),
    .INIT_LUTG1(16'b0011101101111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1481|picorv32_core/reg5_b15_placeOpt_3  (
    .a({_al_u1088_o,_al_u1089_o}),
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,mem_rdata[31]}),
    .c({_al_u1470_o,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u1469_o,\picorv32_core/mem_la_read }),
    .e({\picorv32_core/mem_16bit_buffer [15],\picorv32_core/mem_16bit_buffer [15]}),
    .f({_al_u1481_o_placeOpt_3,open_n6407}));  // ../src/picorv32.v(605)
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTF1("~(~0*~((D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))*~(B)+~0*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*~(B)+~(~0)*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*B+~0*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*B)"),
    //.LUTG0("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTG1("~(~1*~((D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))*~(B)+~1*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*~(B)+~(~1)*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*B+~1*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010011000000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1110111011001111),
    .INIT_LUTG1(16'b0011101101111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1481|picorv32_core/reg5_b15_placeOpt_4  (
    .a({_al_u1088_o,_al_u1089_o}),
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,mem_rdata[31]}),
    .c({_al_u1470_o,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u1469_o,\picorv32_core/mem_la_read }),
    .e({\picorv32_core/mem_16bit_buffer [15],\picorv32_core/mem_16bit_buffer [15]}),
    .f({_al_u1481_o_placeOpt_4,open_n6428}));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUT1("~(~1*~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*~(B)+~1*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)+~(~1)*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B+~1*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B)"),
    .INIT_LUT0(16'b0000001010001010),
    .INIT_LUT1(16'b0011011110111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1485 (
    .a({_al_u1088_o,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,_al_u1088_o}),
    .c({_al_u1439_o,_al_u1439_o}),
    .d({_al_u1440_o,_al_u1440_o}),
    .mi({open_n6446,\picorv32_core/mem_16bit_buffer [13]}),
    .fx({open_n6451,_al_u1485_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))*~(C)+~0*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*~(C)+~(~0)*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*C+~0*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*C)"),
    //.LUT1("~(~1*~((D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))*~(C)+~1*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*~(C)+~(~1)*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*C+~1*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)*C)"),
    .INIT_LUT0(16'b0100000001110000),
    .INIT_LUT1(16'b0100111101111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1485_placeOpt_1 (
    .a({_al_u1440_o,_al_u1440_o}),
    .b({_al_u1088_o,_al_u1088_o}),
    .c({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .d({_al_u1439_o,_al_u1439_o}),
    .mi({open_n6466,\picorv32_core/mem_16bit_buffer [13]}),
    .fx({open_n6471,_al_u1485_o_placeOpt_1}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUT1("~(~1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    .INIT_LUT0(16'b0000001010001010),
    .INIT_LUT1(16'b0101011111011111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1485_placeOpt_2 (
    .a({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({_al_u1088_o,_al_u1088_o}),
    .c({_al_u1439_o,_al_u1439_o}),
    .d({_al_u1440_o,_al_u1440_o}),
    .mi({open_n6486,\picorv32_core/mem_16bit_buffer [13]}),
    .fx({open_n6491,_al_u1485_o_placeOpt_2}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUT1("~(~1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(~1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+~1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    .INIT_LUT0(16'b0000001010001010),
    .INIT_LUT1(16'b0101011111011111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1485_placeOpt_3 (
    .a({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({_al_u1088_o,_al_u1088_o}),
    .c({_al_u1439_o,_al_u1439_o}),
    .d({_al_u1440_o,_al_u1440_o}),
    .mi({open_n6506,\picorv32_core/mem_16bit_buffer [13]}),
    .fx({open_n6511,_al_u1485_o_placeOpt_3}));
  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~C*~(B*D))"),
    //.LUT1("(~B*~C*~A*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110111110101),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1494|picorv32_core/mem_valid_reg  (
    .a({_al_u1493_o,_al_u1557_o}),
    .b({\picorv32_core/mem_state [1],\picorv32_core/mux59_sel_is_5_o }),
    .c({\picorv32_core/mem_state [0],\picorv32_core/n25 }),
    .clk(clk_pad),
    .d({_al_u1089_o,\picorv32_core/mem_la_read }),
    .sr(\picorv32_core/n111 ),
    .f({\picorv32_core/n25 ,open_n6527}),
    .q({open_n6531,\picorv32_core/mem_valid }));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~D))"),
    //.LUT1("(B*~(C*~A))"),
    .INIT_LUT0(16'b1100110000001100),
    .INIT_LUT1(16'b1000110010001100),
    .MODE("LOGIC"))
    \_al_u1496|_al_u1537  (
    .a({_al_u1261_o,open_n6532}),
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .c({_al_u1088_o,_al_u1088_o}),
    .d({open_n6535,_al_u1432_o}),
    .f({_al_u1496_o,_al_u1537_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)"),
    //.LUTF1("D*~A*~C*~B+D*A*~C*~B+D*~A*C*~B+D*A*C*~B"),
    //.LUTG0("(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)"),
    //.LUTG1("D*~A*~C*~B+D*A*~C*~B+D*~A*C*~B+D*A*C*~B+~D*~A*~C*B+D*~A*~C*B+~D*A*~C*B+D*A*~C*B+~D*~A*C*B+D*~A*C*B+~D*A*C*B+D*A*C*B"),
    .INIT_LUTF0(16'b1101110110001000),
    .INIT_LUTF1(16'b0011001100000000),
    .INIT_LUTG0(16'b1101110110001000),
    .INIT_LUTG1(16'b1111111111001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1501|_al_u1519  (
    .a({open_n6554,uart_sel_lutinv_placeOpt_1}),
    .b({uart_sel_lutinv_placeOpt_1,uart_do[30]}),
    .d({memory_out[25],memory_out[30]}),
    .e({uart_do[25],open_n6559}),
    .f({mem_rdata[25],mem_rdata[30]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*D*~C*~B+A*D*~C*~B+~A*D*C*~B+A*D*C*~B+~A*D*~C*B+A*D*~C*B+~A*D*C*B+A*D*C*B"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1505|_al_u1530  (
    .b({uart_do[23],open_n6582}),
    .c({memory_out[23],uart_do[16]}),
    .d({uart_sel_lutinv_placeOpt_3,memory_out[16]}),
    .e({open_n6585,uart_sel_lutinv_placeOpt_3}),
    .f({mem_rdata[23],mem_rdata[16]}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*C*~D+A*B*C*~D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~B*A*~C*~D+B*A*~C*~D+~B*A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~B*A*~C*~D+B*A*~C*~D+~B*A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    .INIT_LUTF0(16'b1010000010100000),
    .INIT_LUTF1(16'b1111101000001010),
    .INIT_LUTG0(16'b1111010111110101),
    .INIT_LUTG1(16'b1111101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1507|_al_u1511  (
    .a({memory_out[22],uart_sel_lutinv_placeOpt_1}),
    .c({uart_sel_lutinv_placeOpt_1,uart_do[20]}),
    .d({uart_do[22],open_n6610}),
    .e({open_n6611,memory_out[20]}),
    .f({mem_rdata[22],mem_rdata[20]}));
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(~0*~B*~C*A))"),
    //.LUTF1("0"),
    //.LUTG0("~(~D*~(~1*~B*~C*A))"),
    //.LUTG1("~A*~D*~B*C+~A*D*~B*C+~A*~D*B*C+~A*D*B*C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100000010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b0101000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1533|picorv32_core/is_beq_bne_blt_bge_bltu_bgeu_reg  (
    .a({\picorv32_core/mem_rdata_latched [4],_al_u1533_o}),
    .b({open_n6632,\picorv32_core/mem_rdata_latched [3]}),
    .c({\picorv32_core/mem_rdata_latched [6],\picorv32_core/n180 }),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({open_n6633,_al_u1532_o}),
    .e({\picorv32_core/mem_rdata_latched [5],\picorv32_core/mem_rdata_latched [2]}),
    .sr(resetn_placeOpt_15),
    .f({_al_u1533_o,open_n6648}),
    .q({open_n6652,\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*C*~D)"),
    //.LUT1("(C*D*A)"),
    .INIT_LUT0(16'b0000000001010000),
    .INIT_LUT1(16'b1010000000000000),
    .MODE("LOGIC"))
    \_al_u1535|_al_u2293  (
    .a({\picorv32_core/mem_rdata_latched [2],_al_u1481_o}),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_2 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_2 }),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_4 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .f({_al_u1535_o,_al_u2293_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*D*~C*~B+A*D*~C*~B"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*~C*D+~A*B*~C*D"),
    //.LUTG0("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*~C*B+A*~D*~C*B"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*~C*D+~A*B*~C*D"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0000010100000101),
    .INIT_LUTG0(16'b0000001100001111),
    .INIT_LUTG1(16'b0000010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1538|_al_u1479  (
    .a({\picorv32_core/mux4_b0_sel_is_0_o ,open_n6675}),
    .b({open_n6676,_al_u1282_o}),
    .c({\picorv32_core/mem_16bit_buffer [14],_al_u1089_o}),
    .d({open_n6679,\picorv32_core/mux3_b16_sel_is_0_o }),
    .e({open_n6680,\picorv32_core/mem_rdata_latched_noshuffle [0]}),
    .f({_al_u1538_o,\picorv32_core/mem_rdata_latched [16]}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~A*~(C*~(~0*~B))))"),
    //.LUT1("(D*~(~A*~(C*~(~1*~B))))"),
    .INIT_LUT0(16'b1110101000000000),
    .INIT_LUT1(16'b1111101000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1539 (
    .a({_al_u1538_o,_al_u1538_o}),
    .b({_al_u1431_o,_al_u1431_o}),
    .c({_al_u1537_o,_al_u1537_o}),
    .d({_al_u1485_o,_al_u1485_o}),
    .mi({open_n6713,_al_u1088_o}),
    .fx({open_n6718,\picorv32_core/mux81_sel_is_1_o }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)*A*~(0)+D*~(B)*C*A*~(0)+D*B*C*A*~(0)+D*~(B)*~(C)*~(A)*0+D*~(B)*C*~(A)*0+D*B*C*~(A)*0+D*~(B)*~(C)*A*0+~(D)*~(B)*C*A*0+D*~(B)*C*A*0+~(D)*B*C*A*0+D*B*C*A*0)"),
    //.LUTF1("(D*A)"),
    //.LUTG0("(D*~(B)*~(C)*A*~(1)+D*~(B)*C*A*~(1)+D*B*C*A*~(1)+D*~(B)*~(C)*~(A)*1+D*~(B)*C*~(A)*1+D*B*C*~(A)*1+D*~(B)*~(C)*A*1+~(D)*~(B)*C*A*1+D*~(B)*C*A*1+~(D)*B*C*A*1+D*B*C*A*1)"),
    //.LUTG1("(D*A)"),
    .INIT_LUTF0(16'b1010001000000000),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b1111001110100000),
    .INIT_LUTG1(16'b1010101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1543|_al_u1541  (
    .a({\picorv32_core/n15_lutinv ,\picorv32_core/mem_state [0]}),
    .b({open_n6721,_al_u1186_o}),
    .c({open_n6722,\picorv32_core/mem_do_rinst }),
    .d({resetn_placeOpt_17,\picorv32_core/mem_xfer_placeOpt_1 }),
    .e({open_n6725,\picorv32_core/mem_state [1]}),
    .f({\picorv32_core/n16 ,\picorv32_core/n15_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(0*C*~(A*~(B*D)))"),
    //.LUT1("(1*C*~(A*~(B*D)))"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1101000001010000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1545 (
    .a({_al_u1088_o,_al_u1088_o}),
    .b({\picorv32_core/mem_xfer_placeOpt_4 ,\picorv32_core/mem_xfer_placeOpt_4 }),
    .c({\picorv32_core/n16 ,\picorv32_core/n16 }),
    .d({\picorv32_core/n180 ,\picorv32_core/n180 }),
    .mi({open_n6758,\picorv32_core/mem_do_rinst }),
    .fx({open_n6763,\picorv32_core/n170 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(A*~(C*D))))"),
    //.LUT1("(B*~(1*~(A*~(C*D))))"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1546 (
    .a({\picorv32_core/mem_xfer_placeOpt_3 ,\picorv32_core/mem_xfer_placeOpt_3 }),
    .b({\picorv32_core/n16 ,\picorv32_core/n16 }),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_5 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_5 }),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_2 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_2 }),
    .mi({open_n6778,_al_u1088_o}),
    .fx({open_n6783,_al_u1546_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(A*~(C*D))))"),
    //.LUT1("(B*~(1*~(A*~(C*D))))"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1546_placeOpt_1 (
    .a({\picorv32_core/mem_xfer_placeOpt_3 ,\picorv32_core/mem_xfer_placeOpt_3 }),
    .b({\picorv32_core/n16 ,\picorv32_core/n16 }),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_5 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_5 }),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_2 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_2 }),
    .mi({open_n6798,_al_u1088_o}),
    .fx({open_n6803,_al_u1546_o_placeOpt_1}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(A*~(C*D))))"),
    //.LUT1("(B*~(1*~(A*~(C*D))))"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1546_placeOpt_2 (
    .a({\picorv32_core/mem_xfer_placeOpt_3 ,\picorv32_core/mem_xfer_placeOpt_3 }),
    .b({\picorv32_core/n16 ,\picorv32_core/n16 }),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_5 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_5 }),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_2 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_2 }),
    .mi({open_n6818,_al_u1088_o}),
    .fx({open_n6823,_al_u1546_o_placeOpt_2}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(A*~(C*D))))"),
    //.LUT1("(B*~(1*~(A*~(C*D))))"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1546_placeOpt_3 (
    .a({\picorv32_core/mem_xfer_placeOpt_3 ,\picorv32_core/mem_xfer_placeOpt_3 }),
    .b({\picorv32_core/n16 ,\picorv32_core/n16 }),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_5 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_5 }),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_2 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_2 }),
    .mi({open_n6838,_al_u1088_o}),
    .fx({open_n6843,_al_u1546_o_placeOpt_3}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(A*~(C*D))))"),
    //.LUT1("(B*~(1*~(A*~(C*D))))"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1546_placeOpt_4 (
    .a({\picorv32_core/mem_xfer_placeOpt_3 ,\picorv32_core/mem_xfer_placeOpt_3 }),
    .b({\picorv32_core/n16 ,\picorv32_core/n16 }),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_5 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_5 }),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_2 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_2 }),
    .mi({open_n6858,_al_u1088_o}),
    .fx({open_n6863,_al_u1546_o_placeOpt_4}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(A*~(C*D))))"),
    //.LUT1("(B*~(1*~(A*~(C*D))))"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1546_placeOpt_5 (
    .a({\picorv32_core/mem_xfer_placeOpt_3 ,\picorv32_core/mem_xfer_placeOpt_3 }),
    .b({\picorv32_core/n16 ,\picorv32_core/n16 }),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_5 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_5 }),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_2 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_2 }),
    .mi({open_n6878,_al_u1088_o}),
    .fx({open_n6883,_al_u1546_o_placeOpt_5}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(A*~(C*D))))"),
    //.LUT1("(B*~(1*~(A*~(C*D))))"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1546_placeOpt_6 (
    .a({\picorv32_core/mem_xfer_placeOpt_3 ,\picorv32_core/mem_xfer_placeOpt_3 }),
    .b({\picorv32_core/n16 ,\picorv32_core/n16 }),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_5 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_5 }),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_2 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_2 }),
    .mi({open_n6898,_al_u1088_o}),
    .fx({open_n6903,_al_u1546_o_placeOpt_6}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(A*~(C*D))))"),
    //.LUT1("(B*~(1*~(A*~(C*D))))"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1546_placeOpt_7 (
    .a({\picorv32_core/mem_xfer_placeOpt_3 ,\picorv32_core/mem_xfer_placeOpt_3 }),
    .b({\picorv32_core/n16 ,\picorv32_core/n16 }),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_5 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_5 }),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_2 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_2 }),
    .mi({open_n6918,_al_u1088_o}),
    .fx({open_n6923,_al_u1546_o_placeOpt_7}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(A*~(C*D))))"),
    //.LUT1("(B*~(1*~(A*~(C*D))))"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1546_placeOpt_8 (
    .a({\picorv32_core/mem_xfer_placeOpt_3 ,\picorv32_core/mem_xfer_placeOpt_3 }),
    .b({\picorv32_core/n16 ,\picorv32_core/n16 }),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_5 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_5 }),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_2 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_2 }),
    .mi({open_n6938,_al_u1088_o}),
    .fx({open_n6943,_al_u1546_o_placeOpt_8}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D)*~(B)*~(C)*~(A)*~(0)+D*~(B)*~(C)*~(A)*~(0)+~(D)*B*~(C)*~(A)*~(0)+D*B*~(C)*~(A)*~(0)+~(D)*~(B)*C*~(A)*~(0)+D*~(B)*C*~(A)*~(0)+~(D)*B*C*~(A)*~(0)+D*B*C*~(A)*~(0)+~(D)*~(B)*~(C)*A*~(0)+D*~(B)*~(C)*A*~(0)+~(D)*B*~(C)*A*~(0)+D*B*~(C)*A*~(0)+~(D)*~(B)*C*A*~(0)+D*~(B)*C*A*~(0)+D*~(B)*~(C)*~(A)*0+D*~(B)*C*~(A)*0+D*B*C*~(A)*0+D*~(B)*~(C)*A*0+D*~(B)*C*A*0)"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(~(D)*~(B)*~(C)*~(A)*~(1)+D*~(B)*~(C)*~(A)*~(1)+~(D)*B*~(C)*~(A)*~(1)+D*B*~(C)*~(A)*~(1)+~(D)*~(B)*C*~(A)*~(1)+D*~(B)*C*~(A)*~(1)+~(D)*B*C*~(A)*~(1)+D*B*C*~(A)*~(1)+~(D)*~(B)*~(C)*A*~(1)+D*~(B)*~(C)*A*~(1)+~(D)*B*~(C)*A*~(1)+D*B*~(C)*A*~(1)+~(D)*~(B)*C*A*~(1)+D*~(B)*C*A*~(1)+D*~(B)*~(C)*~(A)*1+D*~(B)*C*~(A)*1+D*B*C*~(A)*1+D*~(B)*~(C)*A*1+D*~(B)*C*A*1)"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0111111101111111),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b0111001100000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1547|_al_u1548  (
    .a({open_n6946,\picorv32_core/mem_do_prefetch_placeOpt_8 }),
    .b({_al_u1184_o,\picorv32_core/n667_lutinv }),
    .c({open_n6947,_al_u1313_o}),
    .d({\picorv32_core/n662 ,_al_u1547_o}),
    .e({\picorv32_core/n666_lutinv ,\picorv32_core/mem_do_rinst }),
    .f({_al_u1547_o,_al_u1548_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b0000101000001010),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1550|picorv32_core/reg18_b9  (
    .a({\picorv32_core/n663 ,\picorv32_core/n502 [9]}),
    .b({open_n6970,\picorv32_core/n504 [9]}),
    .c({\picorv32_core/decoder_trigger ,\picorv32_core/n500 [9]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({open_n6971,\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .f({_al_u1550_o,open_n6986}),
    .q({open_n6990,\picorv32_core/reg_next_pc [9]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A))"),
    //.LUT1("(~A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUT0(16'b1010111100000000),
    .INIT_LUT1(16'b0001000100000101),
    .MODE("LOGIC"))
    \_al_u1551|_al_u1576  (
    .a({\picorv32_core/is_sb_sh_sw ,_al_u1546_o}),
    .b({\picorv32_core/mem_do_rinst ,open_n6991}),
    .c({\picorv32_core/mem_do_prefetch ,\picorv32_core/mem_do_prefetch }),
    .d({\picorv32_core/is_sll_srl_sra ,_al_u1575_o}),
    .f({_al_u1551_o,\picorv32_core/u625_sel_is_2_o }));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*B*C*~(A)*~(0)+~(D)*B*~(C)*A*~(0)+~(D)*B*C*A*~(0)+D*B*C*A*~(0)+D*B*C*~(A)*0+~(D)*~(B)*~(C)*A*0+D*~(B)*~(C)*A*0+~(D)*B*~(C)*A*0+D*B*~(C)*A*0+~(D)*~(B)*C*A*0+D*~(B)*C*A*0+~(D)*B*C*A*0+D*B*C*A*0)"),
    //.LUTF1("0"),
    //.LUTG0("(D*B*C*~(A)*~(1)+~(D)*B*~(C)*A*~(1)+~(D)*B*C*A*~(1)+D*B*C*A*~(1)+D*B*C*~(A)*1+~(D)*~(B)*~(C)*A*1+D*~(B)*~(C)*A*1+~(D)*B*~(C)*A*1+D*B*~(C)*A*1+~(D)*~(B)*C*A*1+D*~(B)*C*A*1+~(D)*B*C*A*1+D*B*C*A*1)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+A*~B*C*~D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000010001000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1110101010101010),
    .INIT_LUTG1(16'b0000000000100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1552|picorv32_core/reg22_b0  (
    .a({_al_u1551_o,resetn_placeOpt_16}),
    .b({\picorv32_core/sel40_b0/or_or_B4_B5_o_or_B6__o_lutinv ,\picorv32_core/n669_lutinv_placeOpt_4 }),
    .c({\picorv32_core/n665_lutinv ,\picorv32_core/mem_do_prefetch_placeOpt_8 }),
    .clk(clk_pad),
    .d({_al_u1550_o,_al_u1546_o}),
    .e({_al_u1548_o,\picorv32_core/sel40_b0/or_or_B4_B5_o_or_B6__o_lutinv }),
    .sr(\picorv32_core/mux164_b0_sel_is_0_o ),
    .f({_al_u1552_o,open_n7027}),
    .q({open_n7031,\picorv32_core/cpu_state [0]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(B*~(~D*C)))"),
    //.LUT1("(C*~(~A*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111010101110),
    .INIT_LUT1(16'b1111000010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1553|picorv32_core/is_jalr_addi_slti_sltiu_xori_ori_andi_reg  (
    .a({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/instr_jalr }),
    .b({open_n7032,\picorv32_core/is_alu_reg_imm }),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_8 ,\picorv32_core/mem_rdata_q [12]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/is_jalr_addi_slti_sltiu_xori_ori_andi ,\picorv32_core/mem_rdata_q [13]}),
    .f({\picorv32_core/sel23/B2 ,open_n7046}),
    .q({open_n7050,\picorv32_core/is_jalr_addi_slti_sltiu_xori_ori_andi }));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~A*~B*C*~D)"),
    //.LUTF1("~A*~D*~B*~C+A*~D*~B*~C+~A*D*~B*~C+A*D*~B*~C+~A*~D*~B*C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C"),
    //.LUTG0("(~1*~A*~B*C*~D)"),
    //.LUTG1("~A*D*~B*~C+~A*D*~B*C"),
    .INIT_LUTF0(16'b0000000000010000),
    .INIT_LUTF1(16'b0011001100110011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0001000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1554|_al_u1307  (
    .a({\picorv32_core/n524 [7],\picorv32_core/is_lb_lh_lw_lbu_lhu }),
    .b({\picorv32_core/sel23/B2 ,\picorv32_core/is_jalr_addi_slti_sltiu_xori_ori_andi }),
    .c({open_n7051,_al_u1306_o}),
    .d({_al_u1306_o,\picorv32_core/n524 [7]}),
    .e({\picorv32_core/mem_do_rinst ,\picorv32_core/is_lui_auipc_jal }),
    .f({_al_u1554_o,\picorv32_core/n523_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+A*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0)"),
    //.LUT1("(~(A)*~(D)*~(C)*~(B)*~(1)+A*~(D)*~(C)*~(B)*~(1)+~(A)*~(D)*C*~(B)*~(1)+~(A)*~(D)*~(C)*B*~(1)+A*~(D)*~(C)*B*~(1)+~(A)*D*~(C)*B*~(1)+A*D*~(C)*B*~(1)+~(A)*~(D)*C*B*~(1)+A*~(D)*C*B*~(1)+~(A)*D*C*B*~(1)+A*D*C*B*~(1)+~(A)*~(D)*~(C)*~(B)*1+A*~(D)*~(C)*~(B)*1+~(A)*D*~(C)*~(B)*1+A*D*~(C)*~(B)*1+~(A)*~(D)*C*~(B)*1+A*~(D)*C*~(B)*1+~(A)*D*C*~(B)*1+A*D*C*~(B)*1+~(A)*~(D)*~(C)*B*1+A*~(D)*~(C)*B*1+~(A)*D*~(C)*B*1+A*D*~(C)*B*1)"),
    .INIT_LUT0(16'b1111111100010011),
    .INIT_LUT1(16'b0011111100111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1557 (
    .a({_al_u1493_o,_al_u1493_o}),
    .b({\picorv32_core/mem_state [0],\picorv32_core/mem_do_wdata }),
    .c({\picorv32_core/mem_valid ,\picorv32_core/mem_valid }),
    .d({\picorv32_core/mem_do_wdata ,\picorv32_core/mem_state [0]}),
    .mi({open_n7086,\picorv32_core/mem_state [1]}),
    .fx({open_n7091,_al_u1557_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*A*~(0*~(D)*~(B)+0*D*~(B)+~(0)*D*B+0*D*B))"),
    //.LUTF1("(A*D)"),
    //.LUTG0("(C*A*~(1*~(D)*~(B)+1*D*~(B)+~(1)*D*B+1*D*B))"),
    //.LUTG1("(A*D)"),
    .INIT_LUTF0(16'b0010000010100000),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b1010101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1560|_al_u1559  (
    .a({_al_u1559_o,_al_u1481_o}),
    .b({open_n7094,\picorv32_core/mem_rdata_latched$0$_placeOpt_2 }),
    .c({open_n7095,_al_u1483_o_placeOpt_3}),
    .d({_al_u1546_o,\picorv32_core/mem_rdata_latched$1$_placeOpt_3 }),
    .e({open_n7098,_al_u1485_o_placeOpt_1}),
    .f({_al_u1560_o,_al_u1559_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~C*~A))"),
    //.LUT1("~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D)"),
    .INIT_LUT0(16'b1100100011001100),
    .INIT_LUT1(16'b0000111101010101),
    .MODE("LOGIC"))
    \_al_u1563|_al_u1614  (
    .a({\picorv32_core/mem_rdata_q [9],\picorv32_core/mem_xfer_placeOpt_2 }),
    .b({open_n7119,_al_u1613_o}),
    .c({\picorv32_core/mux79_b2/B0_3 ,\picorv32_core/mem_state [0]}),
    .d({\picorv32_core/mem_xfer_placeOpt_2 ,\picorv32_core/mem_state [1]}),
    .f({_al_u1563_o,_al_u1614_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(0*B*A*C))"),
    //.LUT1("(~D*~(1*A*B*C))"),
    .INIT_LUT0(16'b0000000011111111),
    .INIT_LUT1(16'b0000000001111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1565 (
    .a({_al_u1481_o,\picorv32_core/mem_rdata_latched$0$_placeOpt_2 }),
    .b({\picorv32_core/mem_rdata_latched$0$_placeOpt_2 ,_al_u1481_o}),
    .c({\picorv32_core/mem_rdata_latched [4],\picorv32_core/mem_rdata_latched [4]}),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_3 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_3 }),
    .mi({open_n7152,_al_u1483_o_placeOpt_3}),
    .fx({open_n7157,_al_u1565_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(A*B*~(0*~C)))"),
    //.LUTF1("~C*B*~D*~A+~C*B*D*~A+~C*B*~D*A+~C*B*D*A"),
    //.LUTG0("(~D*~(A*B*~(1*~C)))"),
    //.LUTG1("~C*B*~D*~A+~C*B*D*~A"),
    .INIT_LUTF0(16'b0000000001110111),
    .INIT_LUTF1(16'b0000110000001100),
    .INIT_LUTG0(16'b0000000001111111),
    .INIT_LUTG1(16'b0000010000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1567|_al_u1564  (
    .a({\picorv32_core/mem_rdata_latched [6],_al_u1483_o_placeOpt_3}),
    .b({_al_u1565_o,_al_u1481_o}),
    .c({_al_u1564_o,\picorv32_core/mem_rdata_latched$0$_placeOpt_2 }),
    .d({open_n7162,_al_u1563_o}),
    .e({_al_u1566_o,_al_u1485_o_placeOpt_1}),
    .f({_al_u1567_o,_al_u1564_o}));
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~A*~B*~C+D*~A*~B*~C+~D*~A*B*~C+~D*A*B*~C+~D*~A*~B*C+D*~A*~B*C+~D*~A*B*C+~D*A*B*C"),
    //.LUTF1("~B*A*D*~C+B*A*D*~C+~B*A*D*C+B*A*D*C"),
    //.LUTG0("~D*~A*~B*~C+D*~A*~B*~C+~D*~A*~B*C+D*~A*~B*C"),
    //.LUTG1("~B*~A*D*~C+B*~A*D*~C+~B*A*D*~C+B*A*D*~C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001000111011101),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b0001000100010001),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1568|picorv32_core/reg0_b9  (
    .a({_al_u1563_o,_al_u1563_o}),
    .b({open_n7183,_al_u1569_o}),
    .c({\picorv32_core/mux79_b2/B0_3 ,open_n7184}),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_3 ,_al_u1568_o}),
    .e({_al_u1566_o,_al_u1567_o}),
    .f({_al_u1568_o,open_n7201}),
    .q({open_n7205,\picorv32_core/mem_rdata_q [9]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("(~0*C*~(A*~(B*D)))"),
    //.LUT1("(~1*C*~(A*~(B*D)))"),
    .INIT_LUT0(16'b1101000001010000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1569 (
    .a({_al_u1088_o,_al_u1088_o}),
    .b({\picorv32_core/mem_xfer ,\picorv32_core/mem_xfer }),
    .c({\picorv32_core/n16 ,\picorv32_core/n16 }),
    .d({\picorv32_core/n180 ,\picorv32_core/n180 }),
    .mi({open_n7218,_al_u700_o_placeOpt_2}),
    .fx({open_n7223,_al_u1569_o}));
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D)*~(C)*~(A)*~((0*B))+D*~(C)*~(A)*~((0*B))+~(D)*C*~(A)*~((0*B))+~(D)*~(C)*~(A)*(0*B)+D*~(C)*~(A)*(0*B)+~(D)*C*~(A)*(0*B)+D*C*~(A)*(0*B)+D*~(C)*A*(0*B)+D*C*A*(0*B))"),
    //.LUTF1("~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    //.LUTG0("(~(D)*~(C)*~(A)*~((1*B))+D*~(C)*~(A)*~((1*B))+~(D)*C*~(A)*~((1*B))+~(D)*~(C)*~(A)*(1*B)+D*~(C)*~(A)*(1*B)+~(D)*C*~(A)*(1*B)+D*C*~(A)*(1*B)+D*~(C)*A*(1*B)+D*C*A*(1*B))"),
    //.LUTG1("~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010101010101),
    .INIT_LUTF1(16'b0000010111110101),
    .INIT_LUTG0(16'b1100110101010101),
    .INIT_LUTG1(16'b0000010111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1571|picorv32_core/reg0_b8  (
    .a({\picorv32_core/mem_rdata_q [8],_al_u1571_o}),
    .b({open_n7226,_al_u1532_o}),
    .c({\picorv32_core/mem_xfer_placeOpt_2 ,_al_u1559_o}),
    .clk(clk_pad),
    .d({\picorv32_core/mux79_b1/B0_3 ,_al_u1569_o}),
    .e({open_n7228,\picorv32_core/mem_rdata_latched [3]}),
    .f({_al_u1571_o,open_n7244}),
    .q({open_n7248,\picorv32_core/mem_rdata_q [8]}));  // ../src/picorv32.v(508)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*~A))"),
    //.LUT1("~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110001010000),
    .INIT_LUT1(16'b0001000111011101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1573|picorv32_core/reg11_b0  (
    .a({\picorv32_core/mem_rdata_q [7],_al_u803_o}),
    .b({\picorv32_core/mem_xfer_placeOpt_2 ,\picorv32_core/is_sb_sh_sw }),
    .c({open_n7249,\picorv32_core/mem_rdata_q [20]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mux79_b0/B0_3 ,\picorv32_core/mem_rdata_q [7]}),
    .f({_al_u1573_o,open_n7263}),
    .q({open_n7267,\picorv32_core/decoded_imm [0]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~D*~C*~B*~A)"),
    //.LUT1("(1*~D*~C*~B*~A)"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1575 (
    .a({\picorv32_core/n746_lutinv ,\picorv32_core/n746_lutinv }),
    .b({\picorv32_core/n666_lutinv ,\picorv32_core/n666_lutinv }),
    .c({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .d({\picorv32_core/n663 ,\picorv32_core/n663 }),
    .mi({open_n7280,resetn_placeOpt_12}),
    .fx({open_n7285,_al_u1575_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*C*~D))"),
    //.LUT1("(~B*A)"),
    .INIT_LUT0(16'b1100110001001100),
    .INIT_LUT1(16'b0010001000100010),
    .MODE("LOGIC"))
    \_al_u1577|_al_u1578  (
    .a({\picorv32_core/mux59_sel_is_5_o ,resetn_placeOpt_15}),
    .b({\picorv32_core/mem_do_rdata ,_al_u1577_o}),
    .c({open_n7288,\picorv32_core/mem_la_firstword_xfer }),
    .d({open_n7291,\picorv32_core/n180 }),
    .f({_al_u1577_o,\picorv32_core/mux61_sel_is_5_o }));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*~A*~B*C)"),
    //.LUT1("(~1*~D*~A*~B*C)"),
    .INIT_LUT0(16'b0000000000010000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1579 (
    .a({\picorv32_core/mux79_b2/B0_3 ,\picorv32_core/mux79_b2/B0_3 }),
    .b({_al_u1444_o,_al_u1444_o}),
    .c({\picorv32_core/mux79_b1/B0_3 ,\picorv32_core/mux79_b1/B0_3 }),
    .d({\picorv32_core/mux79_b0/B0_3 ,\picorv32_core/mux79_b0/B0_3 }),
    .mi({open_n7322,_al_u1464_o}),
    .fx({open_n7327,_al_u1579_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(0*D*~A*B*~C)"),
    //.LUT1("(1*C*~B*A*~D)"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1580 (
    .a({\picorv32_core/mem_rdata_latched [0],_al_u1481_o}),
    .b({_al_u1481_o,\picorv32_core/mem_rdata_latched [0]}),
    .c({_al_u1483_o,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_4 ,_al_u1483_o}),
    .mi({open_n7342,_al_u1485_o}),
    .fx({open_n7347,_al_u1580_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~A*~C*~B*~D)"),
    //.LUTF1("~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(~1*~A*~C*~B*~D)"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1581|_al_u1605  (
    .a({open_n7350,\picorv32_core/mem_rdata_latched [3]}),
    .b({\picorv32_core/mem_rdata_latched [5],\picorv32_core/mem_rdata_latched [5]}),
    .c({\picorv32_core/mem_rdata_latched [4],\picorv32_core/mem_rdata_latched [4]}),
    .d({\picorv32_core/mem_rdata_latched [6],\picorv32_core/mem_rdata_latched [6]}),
    .e(\picorv32_core/mem_rdata_latched [3:2]),
    .f({_al_u1581_o,_al_u1605_o}));
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0)*~((C*~D*B))+~A*0*~((C*~D*B))+~(~A)*0*(C*~D*B)+~A*0*(C*~D*B))"),
    //.LUTF1("~D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("(~A*~(1)*~((C*~D*B))+~A*1*~((C*~D*B))+~(~A)*1*(C*~D*B)+~A*1*(C*~D*B))"),
    //.LUTG1("~D*~B*~C*~A+~D*~B*C*~A+~D*~B*~C*A+~D*~B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010100010101),
    .INIT_LUTF1(16'b1100110011111111),
    .INIT_LUTG0(16'b0101010111010101),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1583|picorv32_core/reg0_b16  (
    .a({open_n7373,_al_u1583_o}),
    .b({\picorv32_core/mem_xfer ,_al_u1569_o}),
    .c({open_n7374,_al_u1580_o}),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [16],_al_u1579_o}),
    .e({\picorv32_core/mem_rdata_latched [16],\picorv32_core/mem_rdata_latched [6]}),
    .f({_al_u1583_o,open_n7391}),
    .q({open_n7395,\picorv32_core/mem_rdata_q [16]}));  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("D*~B*~C*~A+D*B*~C*~A+D*~B*~C*A+D*B*~C*A"),
    //.LUTF1("~C*~D*~A*~B+~C*D*~A*~B+C*D*~A*~B+~C*~D*A*~B+~C*D*A*~B+C*D*A*~B+~C*~D*~A*B+~C*D*~A*B+C*D*~A*B+~C*~D*A*B+~C*D*A*B+C*D*A*B"),
    //.LUTG0("D*~B*~C*~A+D*~B*~C*A"),
    //.LUTG1("~C*~D*~A*~B+~C*~D*A*~B+~C*~D*~A*B+~C*~D*A*B"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111111100001111),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1585|_al_u2378  (
    .b({open_n7398,_al_u1481_o_placeOpt_1}),
    .c({\picorv32_core/mem_rdata_q [15],_al_u2377_o}),
    .d({\picorv32_core/mem_xfer_placeOpt_2 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_1 }),
    .e({_al_u1481_o_placeOpt_1,_al_u2271_o}),
    .f({_al_u1585_o,_al_u2378_o}));
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0)*~((B*~C*D))+~A*0*~((B*~C*D))+~(~A)*0*(B*~C*D)+~A*0*(B*~C*D))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(~A*~(1)*~((B*~C*D))+~A*1*~((B*~C*D))+~(~A)*1*(B*~C*D)+~A*1*(B*~C*D))"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101010101),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1587|picorv32_core/reg0_b19  (
    .a({\picorv32_core/mem_rdata_latched [19],_al_u1587_o}),
    .b({open_n7421,_al_u1580_o}),
    .c({open_n7422,_al_u1579_o}),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [19],_al_u1569_o}),
    .e({\picorv32_core/mem_xfer_placeOpt_2 ,\picorv32_core/mem_rdata_latched [12]}),
    .f({_al_u1587_o,open_n7439}),
    .q({open_n7443,\picorv32_core/mem_rdata_q [19]}));  // ../src/picorv32.v(508)
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0)*~((B*~C*D))+~A*0*~((B*~C*D))+~(~A)*0*(B*~C*D)+~A*0*(B*~C*D))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(~A*~(1)*~((B*~C*D))+~A*1*~((B*~C*D))+~(~A)*1*(B*~C*D)+~A*1*(B*~C*D))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101010101),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1589|picorv32_core/reg0_b18  (
    .a({open_n7444,_al_u1589_o}),
    .b({open_n7445,_al_u1580_o}),
    .c({\picorv32_core/mem_rdata_latched [18],_al_u1579_o}),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [18],_al_u1569_o}),
    .e({\picorv32_core/mem_xfer_placeOpt_2 ,\picorv32_core/mem_rdata_latched [12]}),
    .f({_al_u1589_o,open_n7462}),
    .q({open_n7466,\picorv32_core/mem_rdata_q [18]}));  // ../src/picorv32.v(508)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A)*~((B*C))+D*A*~((B*C))+~(D)*A*(B*C)+D*A*(B*C))"),
    //.LUT1("~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111110000000),
    .INIT_LUT1(16'b0001000111011101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1591|picorv32_core/reg6_b17  (
    .a({\picorv32_core/mem_rdata_q [17],\picorv32_core/mem_rdata_latched [17]}),
    .b({\picorv32_core/mem_xfer ,\picorv32_core/mem_rdata_latched [0]}),
    .c({open_n7467,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched [17],\picorv32_core/mem_rdata_latched [12]}),
    .f({_al_u1591_o,open_n7481}),
    .q({open_n7485,\picorv32_core/decoded_imm_uj [17]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(0*~B*A*D))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTG0("~(~C*~(1*~B*A*D))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011110000),
    .INIT_LUTF1(16'b0011001100110011),
    .INIT_LUTG0(16'b1111001011110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1594|picorv32_core/is_sb_sh_sw_reg  (
    .a({open_n7486,_al_u1594_o}),
    .b({\picorv32_core/mem_rdata_latched [4],\picorv32_core/mem_rdata_latched [6]}),
    .c({open_n7487,_al_u1566_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({open_n7488,_al_u1593_o}),
    .e({\picorv32_core/mem_rdata_latched [3],\picorv32_core/mem_rdata_latched [5]}),
    .f({_al_u1594_o,open_n7504}),
    .q({open_n7508,\picorv32_core/is_sb_sh_sw }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~A*~D*~B*~C)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u1596|_al_u2403  (
    .a({\picorv32_core/mem_rdata_latched [3],open_n7509}),
    .b({\picorv32_core/mem_rdata_latched [5],_al_u1481_o_placeOpt_3}),
    .c({\picorv32_core/mem_rdata_latched [6],_al_u1483_o_placeOpt_1}),
    .d({\picorv32_core/mem_rdata_latched [4],\picorv32_core/mem_rdata_latched [6]}),
    .f({_al_u1596_o,_al_u2403_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D"),
    //.LUTG0("~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b0101010100001111),
    .INIT_LUTF1(16'b0011000000110000),
    .INIT_LUTG0(16'b0101010100001111),
    .INIT_LUTG1(16'b0011000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1597|_al_u2457  (
    .a({open_n7530,_al_u1483_o_placeOpt_3}),
    .b({_al_u1485_o_placeOpt_1,open_n7531}),
    .c({_al_u1483_o_placeOpt_3,\picorv32_core/mem_rdata_q [14]}),
    .d({open_n7534,\picorv32_core/mem_xfer_placeOpt_2 }),
    .f({_al_u1597_o,_al_u2457_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(C*~(A*~(B*D))))"),
    //.LUTF1("(0*~B*C*~(A*~D))"),
    //.LUTG0("~(1*~(C*~(A*~(B*D))))"),
    //.LUTG1("(1*~B*C*~(A*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1101000001010000),
    .INIT_LUTG1(16'b0011000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1599|picorv32_core/mem_do_rdata_reg  (
    .a({\picorv32_core/mem_do_prefetch ,_al_u1088_o}),
    .b({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_xfer_placeOpt_1 }),
    .c({\picorv32_core/n669_lutinv_placeOpt_4 ,\picorv32_core/n15_lutinv }),
    .ce(\picorv32_core/n747 ),
    .clk(clk_pad),
    .d({_al_u1546_o,\picorv32_core/n180 }),
    .e({resetn_placeOpt_17,resetn_placeOpt_17}),
    .mi({open_n7558,1'b0}),
    .sr(\picorv32_core/n731 ),
    .f({\picorv32_core/n731 ,\picorv32_core/n747 }),
    .q({open_n7573,\picorv32_core/mem_do_rdata }));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~D*~C+~A*B*~D*C"),
    //.LUTF1("(~A*~D*C)"),
    //.LUTG0("~A*~B*~D*~C+~A*B*~D*~C+~A*~B*~D*C+~A*B*~D*C"),
    //.LUTG1("(~A*~D*C)"),
    .INIT_LUTF0(16'b0000000001000100),
    .INIT_LUTF1(16'b0000000001010000),
    .INIT_LUTG0(16'b0000000001010101),
    .INIT_LUTG1(16'b0000000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1601|_al_u2274  (
    .a({_al_u1485_o_placeOpt_3,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .b({open_n7574,_al_u1481_o_placeOpt_2}),
    .c({_al_u1481_o_placeOpt_2,open_n7575}),
    .d({_al_u1483_o_placeOpt_2,_al_u2268_o}),
    .e({open_n7578,_al_u1485_o_placeOpt_3}),
    .f({\picorv32_core/n98_lutinv ,_al_u2274_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+~A*B*C*~D"),
    //.LUTF1("~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*B*~C*~D+~A*B*C*~D"),
    //.LUTG1("~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000000001000100),
    .INIT_LUTF1(16'b1100110000000000),
    .INIT_LUTG0(16'b0000000001000100),
    .INIT_LUTG1(16'b1100110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1602|_al_u2422  (
    .a({open_n7599,_al_u1485_o}),
    .b({_al_u1464_o,_al_u1464_o}),
    .d({_al_u1444_o,_al_u1483_o}),
    .f({_al_u1602_o,_al_u2422_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(0*~A*~C*B*D)"),
    //.LUT1("(1*~B*~C*A*D)"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000001000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1603 (
    .a({_al_u1602_o,\picorv32_core/mem_rdata_latched$1$_placeOpt_3 }),
    .b({\picorv32_core/mem_rdata_latched$1$_placeOpt_3 ,_al_u1602_o}),
    .c({\picorv32_core/mem_rdata_latched [12],\picorv32_core/mem_rdata_latched [12]}),
    .d({\picorv32_core/n98_lutinv ,\picorv32_core/n98_lutinv }),
    .mi({open_n7638,\picorv32_core/mem_rdata_latched$0$_placeOpt_2 }),
    .fx({open_n7643,_al_u1603_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("B*C*~D*~A+~B*~C*D*~A+B*~C*D*~A+~B*C*D*~A+B*C*D*~A+B*C*~D*A+~B*~C*D*A+B*~C*D*A+~B*C*D*A+B*C*D*A"),
    //.LUTF1("~A*~B*~C*D+~A*B*~C*D"),
    //.LUTG0("B*C*~D*~A+B*C*D*~A+B*C*~D*A+B*C*D*A"),
    //.LUTG1("~A*~B*~C*D+~A*B*~C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b0000010100000000),
    .INIT_LUTG0(16'b1100000011000000),
    .INIT_LUTG1(16'b0000010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1604|picorv32_core/instr_lui_reg  (
    .a({\picorv32_core/n180 ,open_n7646}),
    .b({open_n7647,_al_u1535_o}),
    .c({\picorv32_core/mem_rdata_latched [2],_al_u1581_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u1581_o,_al_u1580_o}),
    .e({open_n7648,_al_u1579_o}),
    .f({_al_u1604_o,open_n7664}),
    .q({open_n7668,\picorv32_core/instr_lui }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B*~(D*~(~0*C)))"),
    //.LUT1("(~A*~C*~(D*~(~1*B)))"),
    .INIT_LUT0(16'b0001000000010001),
    .INIT_LUT1(16'b0000000000000101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1606 (
    .a({_al_u1296_o,_al_u1296_o}),
    .b({\picorv32_core/mem_rdata_latched_noshuffle [1],\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_3 ,\picorv32_core/mem_rdata_latched_noshuffle [1]}),
    .d({_al_u1295_o,_al_u1295_o}),
    .mi({open_n7681,_al_u1088_o}),
    .fx({open_n7686,_al_u1606_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~A*~B*~D+~C*A*~B*~D+~C*~A*~B*D+~C*A*~B*D+~C*~A*B*D+~C*A*B*D"),
    //.LUTF1("(~C*~(B*~A))"),
    //.LUTG0("0"),
    //.LUTG1("(~C*~(B*~A))"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b0000101100001011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000101100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1608|_al_u2258  (
    .a({_al_u1546_o,open_n7689}),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_8 ,\picorv32_core/mem_do_prefetch_placeOpt_8 }),
    .c({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_rdata }),
    .d({open_n7692,_al_u1546_o}),
    .e({open_n7693,\picorv32_core/n576 [0]}),
    .f({\picorv32_core/mux132_b0_sel_is_3_o ,_al_u2258_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D))"),
    //.LUT1("(~1*(~(A)*~(D)*~(C)*~(B)+A*~(D)*~(C)*~(B)+~(A)*~(D)*C*~(B)+A*~(D)*C*~(B)+~(A)*D*C*~(B)+A*D*C*~(B)+~(A)*~(D)*~(C)*B+A*~(D)*~(C)*B+~(A)*D*~(C)*B+A*D*~(C)*B+A*~(D)*C*B+A*D*C*B))"),
    .INIT_LUT0(16'b1010111111110011),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1613 (
    .a({\picorv32_core/mem_do_rinst ,\picorv32_core/mem_do_rinst }),
    .b({\picorv32_core/mem_state [1],\picorv32_core/mem_do_wdata }),
    .c({\picorv32_core/mem_state [0],\picorv32_core/mem_state [0]}),
    .d({\picorv32_core/mem_do_wdata ,\picorv32_core/mem_state [1]}),
    .mi({open_n7726,trap_pad}),
    .fx({open_n7731,_al_u1613_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~((A*~D))*~(C)+~(0*~B)*(A*~D)*~(C)+~(~(0*~B))*(A*~D)*C+~(0*~B)*(A*~D)*C)"),
    //.LUTF1("D*C*A*~B+D*C*A*B"),
    //.LUTG0("(~(1*~B)*~((A*~D))*~(C)+~(1*~B)*(A*~D)*~(C)+~(~(1*~B))*(A*~D)*C+~(1*~B)*(A*~D)*C)"),
    //.LUTG1("D*~C*A*~B+D*C*A*~B+D*~C*A*B+D*C*A*B"),
    .INIT_LUTF0(16'b0000111110101111),
    .INIT_LUTF1(16'b1010000000000000),
    .INIT_LUTG0(16'b0000110010101100),
    .INIT_LUTG1(16'b1010101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1617|_al_u1619  (
    .a({\picorv32_core/mem_state [0],_al_u1617_o}),
    .b({open_n7734,\picorv32_core/mem_do_rinst }),
    .c({\picorv32_core/mem_do_rdata ,_al_u1618_o}),
    .d({\picorv32_core/mem_xfer_placeOpt_1 ,\picorv32_core/mem_la_read }),
    .e({\picorv32_core/mem_do_rinst ,\picorv32_core/mem_state [0]}),
    .f({_al_u1617_o,_al_u1619_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(~B*~(~C*~(~D*~A)))"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b0011000000110001),
    .MODE("LOGIC"))
    \_al_u1618|_al_u1128  (
    .a({_al_u1493_o,\picorv32_core/mem_do_wdata }),
    .b(\picorv32_core/mem_state ),
    .c({\picorv32_core/mem_state [0],\picorv32_core/mem_state [1]}),
    .d({\picorv32_core/mem_do_wdata ,resetn_placeOpt_13}),
    .f({_al_u1618_o,_al_u1128_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    //.LUT1("(A*B*~D)"),
    .INIT_LUT0(16'b0001000111011101),
    .INIT_LUT1(16'b0000000010001000),
    .MODE("LOGIC"))
    \_al_u1621|_al_u2465  (
    .a({_al_u1464_o,\picorv32_core/mem_rdata_q [12]}),
    .b({_al_u1444_o,\picorv32_core/mem_xfer_placeOpt_2 }),
    .d({\picorv32_core/mem_rdata_latched [12],\picorv32_core/mem_rdata_latched [12]}),
    .f({_al_u1621_o,_al_u2465_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*C*~D"),
    //.LUTF1("A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTG0("A*~B*C*~D"),
    //.LUTG1("A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b0000111100001110),
    .INIT_LUTG0(16'b0000000000100000),
    .INIT_LUTG1(16'b0000111100001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1622|_al_u1566  (
    .a({_al_u1621_o,_al_u1483_o}),
    .b({\picorv32_core/mem_rdata_latched [5],\picorv32_core/mem_rdata_latched [0]}),
    .c({\picorv32_core/mem_rdata_latched$1$_placeOpt_4 ,_al_u1481_o_placeOpt_4}),
    .d({_al_u1566_o,_al_u1485_o}),
    .f({_al_u1622_o,_al_u1566_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*(D*C*~(A)+~(D)*~(C)*A+D*~(C)*A))"),
    //.LUT1("(~1*A*(D*B*~(C)+~(D)*~(B)*C+D*~(B)*C))"),
    .INIT_LUT0(16'b0100100000001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1623 (
    .a({_al_u1481_o_placeOpt_4,_al_u1483_o}),
    .b({\picorv32_core/mem_rdata_latched [0],_al_u1481_o_placeOpt_4}),
    .c({_al_u1483_o,\picorv32_core/mem_rdata_latched [0]}),
    .d({_al_u1621_o,_al_u1621_o}),
    .mi({open_n7835,_al_u1485_o}),
    .fx({open_n7840,_al_u1623_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D)*~(B)*~(C)*~(A)*~(0)+D*~(B)*~(C)*~(A)*~(0)+~(D)*B*~(C)*~(A)*~(0)+D*B*~(C)*~(A)*~(0)+~(D)*~(B)*~(C)*A*~(0)+D*~(B)*~(C)*A*~(0)+~(D)*B*~(C)*A*~(0)+D*B*~(C)*A*~(0)+~(D)*~(B)*~(C)*~(A)*0+D*~(B)*~(C)*~(A)*0+~(D)*B*~(C)*~(A)*0+D*B*~(C)*~(A)*0+~(D)*~(B)*C*~(A)*0+D*~(B)*C*~(A)*0+~(D)*B*C*~(A)*0+D*B*C*~(A)*0+~(D)*~(B)*~(C)*A*0+D*~(B)*~(C)*A*0+~(D)*B*~(C)*A*0+D*~(B)*C*A*0)"),
    //.LUTF1("0"),
    //.LUTG0("(~(D)*~(B)*~(C)*~(A)*~(1)+D*~(B)*~(C)*~(A)*~(1)+~(D)*B*~(C)*~(A)*~(1)+D*B*~(C)*~(A)*~(1)+~(D)*~(B)*~(C)*A*~(1)+D*~(B)*~(C)*A*~(1)+~(D)*B*~(C)*A*~(1)+D*B*~(C)*A*~(1)+~(D)*~(B)*~(C)*~(A)*1+D*~(B)*~(C)*~(A)*1+~(D)*B*~(C)*~(A)*1+D*B*~(C)*~(A)*1+~(D)*~(B)*C*~(A)*1+D*~(B)*C*~(A)*1+~(D)*B*C*~(A)*1+D*B*C*~(A)*1+~(D)*~(B)*~(C)*A*1+D*~(B)*~(C)*A*1+~(D)*B*~(C)*A*1+D*~(B)*C*A*1)"),
    //.LUTG1("~B*~A*~C*~D+~B*A*~C*~D+~B*~A*C*~D+~B*A*C*~D+~B*~A*~C*D+~B*A*~C*D+~B*~A*C*D+~B*A*C*D"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0111011101011111),
    .INIT_LUTG1(16'b0011001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1624|_al_u2408  (
    .a({open_n7843,_al_u1483_o_placeOpt_2}),
    .b({_al_u1485_o_placeOpt_2,\picorv32_core/mem_rdata_latched [5]}),
    .c({open_n7844,\picorv32_core/mem_rdata_latched [12]}),
    .d({open_n7847,_al_u1579_o}),
    .e({\picorv32_core/mem_rdata_latched [5],_al_u1485_o_placeOpt_2}),
    .f({\picorv32_core/sel10_b3/B1_1 ,_al_u2408_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~C*B*~D*A)"),
    //.LUT1("(~1*~C*B*~D*A)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1627 (
    .a({\picorv32_core/mem_rdata_latched$0$_placeOpt_4 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .b({_al_u1481_o_placeOpt_4,_al_u1481_o_placeOpt_4}),
    .c({_al_u1483_o,_al_u1483_o}),
    .d({_al_u1464_o,_al_u1464_o}),
    .mi({open_n7880,_al_u1485_o}),
    .fx({open_n7885,_al_u1627_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~A*~(C*~(~0*B))))"),
    //.LUTF1("(~A*D*~(C*~(~0*B)))"),
    //.LUTG0("(~D*~(~A*~(C*~(~1*B))))"),
    //.LUTG1("(~A*D*~(C*~(~1*B)))"),
    .INIT_LUTF0(16'b0000000010111010),
    .INIT_LUTF1(16'b0100010100000000),
    .INIT_LUTG0(16'b0000000011111010),
    .INIT_LUTG1(16'b0000010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1632|_al_u1498  (
    .a({_al_u1497_o,_al_u1497_o}),
    .b({\picorv32_core/mem_rdata_latched_noshuffle [5],\picorv32_core/mem_rdata_latched_noshuffle [5]}),
    .c({_al_u1496_o,_al_u1496_o}),
    .d({\picorv32_core/mem_rdata_latched [6],\picorv32_core/mem_rdata_latched [6]}),
    .e({_al_u1088_o,_al_u1088_o}),
    .f({\picorv32_core/n68 [0],_al_u1498_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(0*B*A*~D))"),
    //.LUTF1("(0*~A*~B*C*~D)"),
    //.LUTG0("~(~C*~(1*B*A*~D))"),
    //.LUTG1("(1*~A*~B*C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000011111000),
    .INIT_LUTG1(16'b0000000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1633|picorv32_core/instr_jalr_reg  (
    .a({\picorv32_core/mem_rdata_latched [3],_al_u1605_o}),
    .b({\picorv32_core/mem_rdata_latched [4],\picorv32_core/n98_lutinv }),
    .c({\picorv32_core/n68 [0],_al_u1633_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/n180 ,_al_u1635_o}),
    .e({\picorv32_core/mem_rdata_latched [2],_al_u1606_o}),
    .f({_al_u1633_o,open_n7925}),
    .q({open_n7929,\picorv32_core/instr_jalr }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D*A)"),
    //.LUT1("(~C*~A)"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"))
    \_al_u1634|_al_u2362  (
    .a({_al_u1464_o,_al_u1444_o}),
    .c({_al_u1444_o,_al_u1485_o_placeOpt_1}),
    .d({open_n7934,_al_u1483_o_placeOpt_3}),
    .f({_al_u1634_o,\picorv32_core/mux79_b3/B1_0 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~B*~C*D*A)"),
    //.LUT1("(~1*~A*~C*D*B)"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1635 (
    .a({\picorv32_core/mux79_b2/B0_3 ,_al_u1634_o}),
    .b({_al_u1634_o,\picorv32_core/mux79_b2/B0_3 }),
    .c({\picorv32_core/mux79_b1/B0_3 ,\picorv32_core/mux79_b1/B0_3 }),
    .d({\picorv32_core/mem_rdata_latched [12],\picorv32_core/mem_rdata_latched [12]}),
    .mi({open_n7965,\picorv32_core/mux79_b0/B0_3 }),
    .fx({open_n7970,_al_u1635_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*((D*~C)*~(0)*~(B)+(D*~C)*0*~(B)+~((D*~C))*0*B+(D*~C)*0*B))"),
    //.LUTF1("(D*~(~A*~(C*~(~0*~B))))"),
    //.LUTG0("(A*((D*~C)*~(1)*~(B)+(D*~C)*1*~(B)+~((D*~C))*1*B+(D*~C)*1*B))"),
    //.LUTG1("(D*~(~A*~(C*~(~1*~B))))"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b1110101000000000),
    .INIT_LUTG0(16'b1000101010001000),
    .INIT_LUTG1(16'b1111101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1639|_al_u1640  (
    .a({_al_u1638_o,\picorv32_core/mem_rdata_latched [1]}),
    .b({_al_u1439_o,\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }),
    .c({_al_u1637_o,_al_u1625_o}),
    .d({\picorv32_core/mem_rdata_latched [4],\picorv32_core/sel10_b2/B1_1 }),
    .e({_al_u1088_o,\picorv32_core/mem_rdata_latched [22]}),
    .f({\picorv32_core/sel10_b2/B1_1 ,_al_u1640_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(~B*~(D*~(~0*~A))))"),
    //.LUTF1("(D*~(~B*~(A*~(~0*~C))))"),
    //.LUTG0("(~C*~(~B*~(D*~(~1*~A))))"),
    //.LUTG1("(D*~(~B*~(A*~(~1*~C))))"),
    .INIT_LUTF0(16'b0000111000001100),
    .INIT_LUTF1(16'b1110110000000000),
    .INIT_LUTG0(16'b0000111100001100),
    .INIT_LUTG1(16'b1110111000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1642|_al_u2291  (
    .a({_al_u1637_o,_al_u1439_o}),
    .b({_al_u1638_o,_al_u1638_o}),
    .c({_al_u1439_o,_al_u1481_o_placeOpt_4}),
    .d({\picorv32_core/mem_rdata_latched [3],_al_u1637_o}),
    .e({_al_u1088_o,_al_u1088_o}),
    .f({\picorv32_core/sel10_b1/B1_1 ,_al_u2291_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*((D*~B)*~(0)*~(A)+(D*~B)*0*~(A)+~((D*~B))*0*A+(D*~B)*0*A))"),
    //.LUT1("(B*((D*~C)*~(1)*~(A)+(D*~C)*1*~(A)+~((D*~C))*1*A+(D*~C)*1*A))"),
    .INIT_LUT0(16'b0001000000000000),
    .INIT_LUT1(16'b1000110010001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1643 (
    .a({\picorv32_core/mem_rdata_latched$0$_placeOpt_3 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }),
    .b({\picorv32_core/mem_rdata_latched [1],_al_u1625_o}),
    .c({_al_u1625_o,\picorv32_core/mem_rdata_latched [1]}),
    .d({\picorv32_core/sel10_b1/B1_1 ,\picorv32_core/sel10_b1/B1_1 }),
    .mi({open_n8029,\picorv32_core/mem_rdata_latched [21]}),
    .fx({open_n8034,_al_u1643_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((D*~C)*~(0)*~(B)+(D*~C)*0*~(B)+~((D*~C))*0*B+(D*~C)*0*B))"),
    //.LUT1("(C*((D*~A)*~(1)*~(B)+(D*~A)*1*~(B)+~((D*~A))*1*B+(D*~A)*1*B))"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b1101000011000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1646 (
    .a({_al_u1625_o,\picorv32_core/mem_rdata_latched [1]}),
    .b({\picorv32_core/mem_rdata_latched$0$_placeOpt_3 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }),
    .c({\picorv32_core/mem_rdata_latched [1],_al_u1625_o}),
    .d({\picorv32_core/sel10_b0/B1_1 ,\picorv32_core/sel10_b0/B1_1 }),
    .mi({open_n8049,\picorv32_core/mem_rdata_latched [20]}),
    .fx({open_n8054,_al_u1646_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(~(C)*~(B)*~(A)*~(0)+C*~(B)*~(A)*~(0)+~(C)*B*~(A)*~(0)+C*B*~(A)*~(0)+~(C)*B*A*~(0)+~(C)*B*~(A)*0+C*B*~(A)*0))"),
    //.LUTF1("~C*~B*~D*~A+C*~B*~D*~A+~C*B*~D*~A+C*B*~D*~A+~C*~B*D*~A+C*~B*D*~A+~C*B*D*~A+C*B*D*~A+~C*~B*~D*A+C*~B*~D*A+~C*~B*D*A+C*~B*D*A"),
    //.LUTG0("(D*(~(C)*~(B)*~(A)*~(1)+C*~(B)*~(A)*~(1)+~(C)*B*~(A)*~(1)+C*B*~(A)*~(1)+~(C)*B*A*~(1)+~(C)*B*~(A)*1+C*B*~(A)*1))"),
    //.LUTG1("~C*~B*D*~A+C*~B*D*~A+~C*B*D*~A+C*B*D*~A+~C*~B*D*A+C*~B*D*A"),
    .INIT_LUTF0(16'b0101110100000000),
    .INIT_LUTF1(16'b0111011101110111),
    .INIT_LUTG0(16'b0100010000000000),
    .INIT_LUTG1(16'b0111011100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1648|_al_u1649  (
    .a({\picorv32_core/mem_rdata_latched$1$_placeOpt_3 ,_al_u1481_o}),
    .b({\picorv32_core/mem_rdata_latched$0$_placeOpt_2 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_2 }),
    .c({open_n8057,_al_u1602_o}),
    .d({_al_u1483_o_placeOpt_3,_al_u1648_o}),
    .e({_al_u1485_o_placeOpt_1,_al_u1483_o_placeOpt_3}),
    .f({_al_u1648_o,_al_u1649_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B)"),
    //.LUT1("(~B*D*A)"),
    .INIT_LUT0(16'b0000001100000011),
    .INIT_LUT1(16'b0010001000000000),
    .MODE("LOGIC"))
    \_al_u1651|_al_u1650  (
    .a({_al_u1650_o,open_n8080}),
    .b({\picorv32_core/mem_rdata_latched [12],\picorv32_core/mem_rdata_latched$1$_placeOpt_3 }),
    .c({open_n8081,\picorv32_core/mem_rdata_latched$0$_placeOpt_1 }),
    .d({_al_u1498_o,open_n8084}),
    .f({_al_u1651_o,_al_u1650_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~B*A*C*~D)"),
    //.LUT1("(~1*~B*A*C*~D)"),
    .INIT_LUT0(16'b0000000000100000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1652 (
    .a({\picorv32_core/mem_rdata_latched [4],\picorv32_core/mem_rdata_latched [4]}),
    .b({\picorv32_core/mem_rdata_latched [3],\picorv32_core/mem_rdata_latched [3]}),
    .c({_al_u1498_o,_al_u1498_o}),
    .d({\picorv32_core/n180 ,\picorv32_core/n180 }),
    .mi({open_n8115,\picorv32_core/mem_rdata_latched [2]}),
    .fx({open_n8120,_al_u1652_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(~D*~B*C*A))"),
    //.LUT1("(1*~(~D*~B*C*A))"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1111111111011111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1653 (
    .a({_al_u1634_o,_al_u1634_o}),
    .b({\picorv32_core/mux79_b2/B0_3 ,\picorv32_core/mux79_b2/B0_3 }),
    .c({\picorv32_core/mux79_b1/B0_3 ,\picorv32_core/mux79_b1/B0_3 }),
    .d({\picorv32_core/mux79_b0/B0_3 ,\picorv32_core/mux79_b0/B0_3 }),
    .mi({open_n8135,_al_u1485_o_placeOpt_1}),
    .fx({open_n8140,_al_u1653_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~C*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D))"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~A*~C*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D))"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b1111000010101010),
    .INIT_LUTG0(16'b0000010100000100),
    .INIT_LUTG1(16'b1111000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1656|_al_u1712  (
    .a({memory_out[15],\picorv32_core/mem_wordsize [1]}),
    .b({open_n8143,memory_out[15]}),
    .c({uart_do[15],_al_u1663_o}),
    .d({uart_sel_lutinv_placeOpt_1,uart_sel_lutinv_placeOpt_1}),
    .e({open_n8146,uart_do[15]}),
    .f({mem_rdata[15],_al_u1712_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(A*~B)"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0010001000100010),
    .MODE("LOGIC"))
    \_al_u1657|_al_u790  (
    .a({\picorv32_core/mem_wordsize [1],\picorv32_core/mem_wordsize [1]}),
    .b({\picorv32_core/mem_wordsize [0],\picorv32_core/mem_wordsize [0]}),
    .f({_al_u1657_o,\picorv32_core/n734_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)"),
    //.LUT1("(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)"),
    .INIT_LUT0(16'b1111010110100000),
    .INIT_LUT1(16'b1101110110001000),
    .MODE("LOGIC"))
    \_al_u1659|_al_u1813  (
    .a({uart_sel_lutinv_placeOpt_3,uart_sel_lutinv_placeOpt_3}),
    .b({uart_do[7],open_n8191}),
    .c({open_n8192,uart_do[10]}),
    .d({memory_out[7],memory_out[10]}),
    .f({mem_rdata[7],mem_rdata[10]}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*D*~C+A*B*D*~C+A*~B*D*C+A*B*D*C"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    //.LUTG0("~A*~B*~D*~C+~A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+~A*B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b1010101000000000),
    .INIT_LUTF1(16'b0000001100001111),
    .INIT_LUTG0(16'b1111111101010101),
    .INIT_LUTG1(16'b0011001111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1661|_al_u1729  (
    .a({open_n8213,uart_sel_lutinv_placeOpt_3}),
    .b({_al_u1660_o,open_n8214}),
    .c({mem_rdata[7],open_n8215}),
    .d({mem_rdata[23],uart_do[3]}),
    .e({_al_u1136_o,memory_out[3]}),
    .f({_al_u1661_o,mem_rdata[3]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1010101011001100),
    .MODE("LOGIC"))
    \_al_u1662|_al_u1732  (
    .a({uart_do[9],open_n8238}),
    .b({memory_out[9],memory_out[11]}),
    .c({open_n8239,uart_do[11]}),
    .d({uart_sel_lutinv,uart_sel_lutinv}),
    .f({mem_rdata[9],mem_rdata[11]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*A)"),
    //.LUTF1("A*~B*~D*C+A*B*~D*C+A*~B*D*C+A*B*D*C"),
    //.LUTG0("(~B*A)"),
    //.LUTG1("A*~B*~D*C+A*B*~D*C+A*~B*D*C+A*B*D*C"),
    .INIT_LUTF0(16'b0010001000100010),
    .INIT_LUTF1(16'b1010000010100000),
    .INIT_LUTG0(16'b0010001000100010),
    .INIT_LUTG1(16'b1010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1663|_al_u1733  (
    .a({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .b({open_n8260,\picorv32_core/pcpi_rs1$1$ }),
    .c({\picorv32_core/mem_wordsize [0],open_n8261}),
    .f({_al_u1663_o,\picorv32_core/n40 [1]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~1*~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUT0(16'b0011001000010000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1664 (
    .a({\picorv32_core/latched_is_lb ,_al_u1663_o}),
    .b({_al_u1663_o,\picorv32_core/latched_is_lb }),
    .c({mem_rdata[9],mem_rdata[9]}),
    .d({mem_rdata[25],mem_rdata[25]}),
    .mi({open_n8300,\picorv32_core/mem_wordsize [1]}),
    .fx({open_n8305,_al_u1664_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(A*~(C*~D)))"),
    //.LUT1("(~A*~(B*~(C*~D)))"),
    .INIT_LUT0(16'b0001000100110001),
    .INIT_LUT1(16'b0001000101010001),
    .MODE("LOGIC"))
    \_al_u1665|_al_u1877  (
    .a({_al_u1664_o,\picorv32_core/latched_is_lb }),
    .b({\picorv32_core/latched_is_lb ,_al_u1876_o}),
    .c({_al_u1661_o,_al_u1661_o}),
    .d({_al_u1658_o,_al_u1658_o}),
    .f({_al_u1665_o,_al_u1877_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1668|picorv32_core/reg15_b9  (
    .a({_al_u1667_o,_al_u1666_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycle }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [9]}),
    .e({\picorv32_core/pcpi_rs1$9$ ,\picorv32_core/count_instr [41]}),
    .mi({open_n8330,\picorv32_core/n459 [9]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1668_o,_al_u1667_o}),
    .q({open_n8345,\picorv32_core/count_cycle [9]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(A*B))"),
    //.LUTF1("0"),
    //.LUTG0("(C*~(A*B))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b0111000001110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0111000001110000),
    .INIT_LUTG1(16'b0011111100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1669|_al_u1895  (
    .a({open_n8346,\picorv32_core/n543 [1]}),
    .b({\picorv32_core/n666_lutinv ,\picorv32_core/n666_lutinv }),
    .c({\picorv32_core/n543 [9],_al_u1894_o}),
    .e({_al_u1668_o,open_n8351}),
    .f({_al_u1669_o,_al_u1895_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b1111101000001010),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b1111101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1671|_al_u704  (
    .a({memory_out[8],\picorv32_core/n30 [4]}),
    .c({uart_sel_lutinv,\picorv32_core/pcpi_rs1$6$ }),
    .d({uart_do[8],open_n8376}),
    .e({open_n8377,_al_u700_o}),
    .f({mem_rdata[8],mem_la_addr[6]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~1*~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1672 (
    .a({\picorv32_core/latched_is_lb ,\picorv32_core/latched_is_lb }),
    .b({_al_u1663_o,_al_u1663_o}),
    .c({mem_rdata[24],mem_rdata[8]}),
    .d({mem_rdata[8],mem_rdata[24]}),
    .mi({open_n8410,\picorv32_core/mem_wordsize [1]}),
    .fx({open_n8415,_al_u1672_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000001100000011),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1673|picorv32_core/reg13_b8  (
    .a({open_n8418,_al_u1677_o}),
    .b({\picorv32_core/latched_is_lb ,\picorv32_core/n669_lutinv }),
    .c({_al_u1672_o,_al_u1673_o}),
    .clk(clk_pad),
    .d({_al_u1658_o,\picorv32_core/n580 }),
    .e({_al_u1661_o,resetn_placeOpt_10}),
    .f({_al_u1673_o,open_n8435}),
    .q({open_n8439,\picorv32_core/reg_out [8]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1676|picorv32_core/reg15_b40  (
    .a({_al_u1675_o,_al_u1674_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycleh }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [40]}),
    .e({\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/count_instr [8]}),
    .mi({open_n8442,\picorv32_core/n459 [40]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1676_o,_al_u1675_o}),
    .q({open_n8457,\picorv32_core/count_cycle [40]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*A))"),
    //.LUT1("(A*~(C*D))"),
    .INIT_LUT0(16'b0101111100000000),
    .INIT_LUT1(16'b0000101010101010),
    .MODE("LOGIC"))
    \_al_u1677|_al_u1888  (
    .a({_al_u1676_o,\picorv32_core/n666_lutinv }),
    .c({\picorv32_core/n543 [8],\picorv32_core/n543 [10]}),
    .d({\picorv32_core/n666_lutinv ,_al_u1887_o}),
    .f({_al_u1677_o,_al_u1888_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010101010101010),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1679|picorv32_core/reg13_b7  (
    .a({_al_u1661_o,_al_u1683_o}),
    .b({open_n8480,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .c({open_n8481,_al_u1679_o}),
    .clk(clk_pad),
    .d({open_n8483,\picorv32_core/n580 }),
    .e({_al_u1658_o,resetn_placeOpt_12}),
    .f({_al_u1679_o,open_n8499}),
    .q({open_n8503,\picorv32_core/reg_out [7]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1682|picorv32_core/reg15_b7  (
    .a({_al_u1681_o,_al_u1680_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycle }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [7]}),
    .e({\picorv32_core/pcpi_rs1$7$ ,\picorv32_core/count_instr [39]}),
    .mi({open_n8506,\picorv32_core/n459 [7]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1682_o,_al_u1681_o}),
    .q({open_n8521,\picorv32_core/count_cycle [7]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*A))"),
    //.LUT1("(D*~(A*C))"),
    .INIT_LUT0(16'b0101111100000000),
    .INIT_LUT1(16'b0101111100000000),
    .MODE("LOGIC"))
    \_al_u1683|_al_u1881  (
    .a({\picorv32_core/n543 [7],\picorv32_core/n666_lutinv }),
    .c({\picorv32_core/n666_lutinv ,\picorv32_core/n543 [11]}),
    .d({_al_u1682_o,_al_u1880_o}),
    .f({_al_u1683_o,_al_u1881_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D"),
    //.LUTG0("(~1*~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b0000000010101010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111111110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1685|_al_u1855  (
    .a({memory_out[14],\picorv32_core/latched_is_lb }),
    .b({open_n8544,_al_u1663_o}),
    .c({open_n8545,mem_rdata[30]}),
    .d({uart_sel_lutinv_placeOpt_1,mem_rdata[14]}),
    .e({uart_do[14],\picorv32_core/mem_wordsize [1]}),
    .f({mem_rdata[14],_al_u1855_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*B*(D*~(C)*~(0)+D*C*~(0)+~(D)*C*0+D*C*0))"),
    //.LUTF1("(A*B*(D*~(C)*~(0)+D*C*~(0)+~(D)*C*0+D*C*0))"),
    //.LUTG0("(A*B*(D*~(C)*~(1)+D*C*~(1)+~(D)*C*1+D*C*1))"),
    //.LUTG1("(A*B*(D*~(C)*~(1)+D*C*~(1)+~(D)*C*1+D*C*1))"),
    .INIT_LUTF0(16'b1000100000000000),
    .INIT_LUTF1(16'b1000100000000000),
    .INIT_LUTG0(16'b1000000010000000),
    .INIT_LUTG1(16'b1000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1686|_al_u1658  (
    .a({\picorv32_core/pcpi_rs1$0$ ,\picorv32_core/pcpi_rs1$0$ }),
    .b({_al_u1657_o,_al_u1657_o}),
    .c({mem_rdata[30],mem_rdata[31]}),
    .d({mem_rdata[14],mem_rdata[15]}),
    .e({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$1$ }),
    .f({_al_u1686_o,_al_u1658_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~((B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D))*~(C)+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*~(C)+~(A)*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C)"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    //.LUTG0("(A*~((B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D))*~(C)+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*~(C)+~(A)*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C)"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b0000101011001010),
    .INIT_LUTF1(16'b0010001000110000),
    .INIT_LUTG0(16'b1111101011001010),
    .INIT_LUTG1(16'b0010001000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1687|_al_u1256  (
    .a({uart_do[6],\picorv32_core/mem_rdata_q [6]}),
    .b({_al_u1136_o,memory_out[6]}),
    .c({memory_out[6],\picorv32_core/mem_xfer_placeOpt_1 }),
    .d({uart_sel_lutinv_placeOpt_1,uart_sel_lutinv_placeOpt_1}),
    .e({open_n8592,uart_do[6]}),
    .f({_al_u1687_o,\picorv32_core/mem_rdata_latched_noshuffle [6]}));
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D"),
    //.LUTG0("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010011000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1110111011001111),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1688|picorv32_core/reg5_b6  (
    .a({open_n8613,_al_u1089_o}),
    .b({mem_rdata[22],mem_rdata[22]}),
    .c({_al_u1687_o,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u1686_o,\picorv32_core/mem_la_read }),
    .e({_al_u1660_o,\picorv32_core/mem_16bit_buffer [6]}),
    .f({_al_u1688_o,open_n8629}),
    .q({open_n8633,\picorv32_core/mem_16bit_buffer [6]}));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(~(0*C*B)*~(D*A))"),
    //.LUT1("(~(1*C*B)*~(D*A))"),
    .INIT_LUT0(16'b0101010111111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1689 (
    .a({\picorv32_core/n666_lutinv ,\picorv32_core/n666_lutinv }),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .c({_al_u1313_o,_al_u1313_o}),
    .d({\picorv32_core/n543 [6],\picorv32_core/n543 [6]}),
    .mi({open_n8646,\picorv32_core/pcpi_rs1$6$ }),
    .fx({open_n8651,_al_u1689_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("0"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b1111111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1692|picorv32_core/reg15_b38  (
    .a({open_n8654,_al_u1690_o}),
    .b({open_n8655,\picorv32_core/instr_rdcycleh }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1691_o,\picorv32_core/count_cycle [38]}),
    .e({_al_u1689_o,\picorv32_core/count_instr [6]}),
    .mi({open_n8658,\picorv32_core/n459 [38]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1692_o,_al_u1691_o}),
    .q({open_n8673,\picorv32_core/count_cycle [38]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~C*B*~D+A*C*B*~D+A*~C*B*D+A*C*B*D"),
    //.LUTF1("A*B*~C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG1("A*B*~C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b1101110110001000),
    .INIT_LUTG0(16'b1101110111011101),
    .INIT_LUTG1(16'b1101110110001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1694|_al_u1703  (
    .a({uart_sel_lutinv_placeOpt_1,uart_sel_lutinv_placeOpt_1}),
    .b(uart_do[13:12]),
    .d({memory_out[13],open_n8678}),
    .e({open_n8679,memory_out[12]}),
    .f(mem_rdata[13:12]));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("(A*B*(D*~(C)*~(0)+D*C*~(0)+~(D)*C*0+D*C*0))"),
    //.LUTG0("(~1*~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("(A*B*(D*~(C)*~(1)+D*C*~(1)+~(D)*C*1+D*C*1))"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1000100000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1695|_al_u1862  (
    .a({\picorv32_core/pcpi_rs1$0$ ,\picorv32_core/latched_is_lb }),
    .b({_al_u1657_o,_al_u1663_o}),
    .c({mem_rdata[29],mem_rdata[29]}),
    .d({mem_rdata[13],mem_rdata[13]}),
    .e({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/mem_wordsize [1]}),
    .f({_al_u1695_o,_al_u1862_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~A*~D*~(B*C))"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b0000000000010101),
    .MODE("LOGIC"))
    \_al_u1697|_al_u1696  (
    .a({_al_u1696_o,uart_do[5]}),
    .b({_al_u1660_o,memory_out[5]}),
    .c({mem_rdata[21],_al_u1136_o}),
    .d({_al_u1695_o,uart_sel_lutinv_placeOpt_1}),
    .f({_al_u1697_o,_al_u1696_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1700|picorv32_core/reg15_b37  (
    .a({_al_u1699_o,_al_u1698_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycleh }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [37]}),
    .e({\picorv32_core/pcpi_rs1$5$ ,\picorv32_core/count_instr [5]}),
    .mi({open_n8744,\picorv32_core/n459 [37]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1700_o,_al_u1699_o}),
    .q({open_n8759,\picorv32_core/count_cycle [37]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*~C*A+B*~D*~C*A+~B*D*~C*A+B*D*~C*A+~B*~D*C*A+B*~D*C*A+~B*D*C*A+B*D*C*A"),
    //.LUTF1("0"),
    //.LUTG0("~B*~D*~C*A+B*~D*~C*A+~B*~D*C*A+B*~D*C*A"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+~A*~D*C*B+A*~D*C*B+~A*D*C*B"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000010101010),
    .INIT_LUTG1(16'b0101010111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1701|_al_u1874  (
    .a({\picorv32_core/n543 [5],_al_u1873_o}),
    .d({\picorv32_core/n666_lutinv ,\picorv32_core/n666_lutinv }),
    .e({_al_u1700_o,\picorv32_core/n543 [12]}),
    .f({_al_u1701_o,_al_u1874_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*B*(C*~(D)*~(0)+C*D*~(0)+~(C)*D*0+C*D*0))"),
    //.LUT1("(A*B*(C*~(D)*~(1)+C*D*~(1)+~(C)*D*1+C*D*1))"),
    .INIT_LUT0(16'b1000000010000000),
    .INIT_LUT1(16'b1000100000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1704 (
    .a({\picorv32_core/pcpi_rs1$0$ ,\picorv32_core/pcpi_rs1$0$ }),
    .b({_al_u1657_o,_al_u1657_o}),
    .c({mem_rdata[12],mem_rdata[12]}),
    .d({mem_rdata[28],mem_rdata[28]}),
    .mi({open_n8798,\picorv32_core/pcpi_rs1$1$ }),
    .fx({open_n8803,_al_u1704_o}));
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(~B)"),
    //.LUT1("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001100110011),
    .INIT_LUT1(16'b0000101000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1705|uart/reg3_b4  (
    .a({uart_do[4],open_n8806}),
    .b({memory_out[4],mem_la_wdata[4]}),
    .c({_al_u1136_o,open_n8807}),
    .ce(\uart/mux15_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({uart_sel_lutinv_placeOpt_1,open_n8808}),
    .mi({open_n8819,mem_la_wdata[4]}),
    .f({_al_u1705_o,n17[4]}),
    .q({open_n8824,\uart/uart_odr [4]}));  // ../src/uart.v(102)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("~C*~A*~D*~B+~C*A*~D*~B+~C*~A*~D*B+~C*A*~D*B"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("~C*~A*~D*~B+~C*A*~D*~B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1706|picorv32_core/reg13_b4  (
    .a({open_n8825,_al_u1710_o}),
    .b({_al_u1660_o,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .c({_al_u1704_o,_al_u1706_o}),
    .clk(clk_pad),
    .d({_al_u1705_o,\picorv32_core/n580 }),
    .e({mem_rdata[20],resetn_placeOpt_13}),
    .f({_al_u1706_o,open_n8842}),
    .q({open_n8846,\picorv32_core/reg_out [4]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1709|picorv32_core/reg15_b4  (
    .a({_al_u1708_o,_al_u1707_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycle }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [4]}),
    .e({\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/count_instr [36]}),
    .mi({open_n8849,\picorv32_core/n459 [4]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1709_o,_al_u1708_o}),
    .q({open_n8864,\picorv32_core/count_cycle [4]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTF1("0"),
    //.LUTG0("~A*~C*~B*D+A*~C*~B*D+~A*~C*B*D+A*~C*B*D"),
    //.LUTG1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*~A*~C*D+B*~A*~C*D+~B*A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0101111101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1710|_al_u1867  (
    .a({\picorv32_core/n666_lutinv ,open_n8865}),
    .c({\picorv32_core/n543 [4],\picorv32_core/n666_lutinv }),
    .d({open_n8870,_al_u1866_o}),
    .e({_al_u1709_o,\picorv32_core/n543 [13]}),
    .f({_al_u1710_o,_al_u1867_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(A*~C*D)"),
    .INIT_LUT0(16'b1100100011101110),
    .INIT_LUT1(16'b0000101000000000),
    .MODE("LOGIC"))
    \_al_u1713|_al_u1140  (
    .a({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/mem_wordsize [0]}),
    .b({open_n8891,\picorv32_core/mem_wordsize [1]}),
    .c({\picorv32_core/mem_wordsize [1],\picorv32_core/pcpi_rs1$0$ }),
    .d({\picorv32_core/mem_wordsize [0],\picorv32_core/pcpi_rs1$1$ }),
    .f({_al_u1713_o,_al_u1140_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+~A*B*C*~D+~A*B*~C*D+~A*B*C*D"),
    //.LUTF1("0"),
    //.LUTG0("A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*D*~B*~C+A*D*~B*~C+A*~D*B*~C+~A*D*B*~C+A*D*B*~C+~A*D*~B*C+A*D*~B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    .INIT_LUTF0(16'b0100010001000100),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1111111110001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1714|_al_u1517  (
    .a({mem_rdata[31],uart_sel_lutinv_placeOpt_1}),
    .b({_al_u1713_o,memory_out[31]}),
    .d({_al_u1712_o,open_n8916}),
    .e({\picorv32_core/latched_is_lh ,uart_do[31]}),
    .f({\picorv32_core/sel27_b16/B1 ,mem_rdata[31]}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("(~B*~D*~(0*~(A*~C)))"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("(~B*~D*~(1*~(A*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1716|picorv32_core/reg13_b31  (
    .a({_al_u1661_o,_al_u1720_o}),
    .b({\picorv32_core/sel27_b31/B2 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .c({_al_u1658_o,_al_u1716_o}),
    .clk(clk_pad),
    .d({\picorv32_core/sel27_b16/B1 ,\picorv32_core/n580 }),
    .e({\picorv32_core/latched_is_lb ,resetn_placeOpt_12}),
    .f({_al_u1716_o,open_n8953}),
    .q({open_n8957,\picorv32_core/reg_out [31]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~D*~B*~C+A*~D*~B*~C+~A*D*~B*~C+A*D*~B*~C+~A*~D*B*~C+~A*D*B*~C+~A*~D*~B*C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C+~A*~D*B*C+~A*D*B*C"),
    //.LUTF1("(~(0*D*B)*~(C*A))"),
    //.LUTG0("~A*~D*~B*~C+A*~D*~B*~C+~A*D*~B*~C+A*D*~B*~C+~A*~D*B*~C+~A*D*B*~C"),
    //.LUTG1("(~(1*D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011101110111),
    .INIT_LUTF1(16'b0101111101011111),
    .INIT_LUTG0(16'b0000011100000111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1717|picorv32_core/reg15_b2  (
    .a({\picorv32_core/n666_lutinv ,\picorv32_core/instr_rdcycle }),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/count_cycle [2]}),
    .c({\picorv32_core/n543 [31],\picorv32_core/count_instr [34]}),
    .clk(clk_pad),
    .d({_al_u1313_o,open_n8959}),
    .e({\picorv32_core/pcpi_rs1$31$ ,\picorv32_core/instr_rdinstrh }),
    .mi({open_n8961,\picorv32_core/n459 [2]}),
    .sr(resetn_placeOpt_8),
    .f({_al_u1717_o,_al_u1815_o}),
    .q({open_n8976,\picorv32_core/count_cycle [2]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(~D*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(~D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010101000001010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b1010101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1720|picorv32_core/reg15_b31  (
    .a({_al_u1717_o,_al_u1718_o}),
    .b({open_n8977,\picorv32_core/instr_rdcycle }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1719_o,\picorv32_core/count_cycle [31]}),
    .e({open_n8979,\picorv32_core/count_instr [63]}),
    .mi({open_n8981,\picorv32_core/n459 [31]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1720_o,_al_u1719_o}),
    .q({open_n8996,\picorv32_core/count_cycle [31]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~B*~(0*~(C*~D)))"),
    //.LUTF1("0"),
    //.LUTG0("(~A*~B*~(1*~(C*~D)))"),
    //.LUTG1("A*B*~C*~D+A*B*C*~D+A*B*~C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0001000100010001),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000010000),
    .INIT_LUTG1(16'b1000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1722|_al_u1723  (
    .a({mem_rdata[30],\picorv32_core/sel27_b30/B2 }),
    .b({\picorv32_core/latched_is_lu ,\picorv32_core/sel27_b16/B1 }),
    .c({open_n8997,_al_u1661_o}),
    .d({open_n9000,_al_u1658_o}),
    .e({\picorv32_core/n734_lutinv ,\picorv32_core/latched_is_lb }),
    .f({\picorv32_core/sel27_b30/B2 ,_al_u1723_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~B*~(0*C)*~(~A*D))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~B*~(1*C)*~(~A*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0010001000110011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1727|picorv32_core/reg15_b30  (
    .a({_al_u1726_o,_al_u1725_o}),
    .b({\picorv32_core/sel43_b30/B2 ,\picorv32_core/instr_rdcycle }),
    .c({\picorv32_core/n666_lutinv ,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({\picorv32_core/n664_lutinv_placeOpt_1 ,\picorv32_core/count_cycle [30]}),
    .e({\picorv32_core/n543 [30],\picorv32_core/count_instr [62]}),
    .mi({open_n9023,\picorv32_core/n459 [30]}),
    .sr(resetn_placeOpt_8),
    .f({_al_u1727_o,_al_u1726_o}),
    .q({open_n9038,\picorv32_core/count_cycle [30]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(~A*D)*~(B*C))"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0010101000111111),
    .MODE("LOGIC"))
    \_al_u1730|_al_u1513  (
    .a({_al_u1136_o,open_n9039}),
    .b({_al_u1660_o,memory_out[19]}),
    .c({mem_rdata[19],uart_do[19]}),
    .d({mem_rdata[3],uart_sel_lutinv_placeOpt_3}),
    .f({_al_u1730_o,mem_rdata[19]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*B*D)"),
    //.LUTF1("(A*B*C)"),
    //.LUTG0("(A*B*D)"),
    //.LUTG1("(A*B*C)"),
    .INIT_LUTF0(16'b1000100000000000),
    .INIT_LUTF1(16'b1000000010000000),
    .INIT_LUTG0(16'b1000100000000000),
    .INIT_LUTG1(16'b1000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1731|_al_u1899  (
    .a({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$1$ }),
    .b({\picorv32_core/pcpi_rs1$0$ ,\picorv32_core/pcpi_rs1$0$ }),
    .c({mem_rdata[27],open_n9060}),
    .d({open_n9063,mem_rdata[24]}),
    .f({_al_u1731_o,_al_u1899_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(0*~(~C*~(A*B))))"),
    //.LUT1("(D*~(1*~(~C*~(A*B))))"),
    .INIT_LUT0(16'b1111111100000000),
    .INIT_LUT1(16'b0000011100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1734 (
    .a({\picorv32_core/n40 [1],\picorv32_core/n40 [1]}),
    .b({mem_rdata[11],mem_rdata[11]}),
    .c({_al_u1731_o,_al_u1731_o}),
    .d({_al_u1730_o,_al_u1730_o}),
    .mi({open_n9098,_al_u1657_o}),
    .fx({open_n9103,_al_u1734_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*C*A)*~(~D*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*C*A)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1111111100110011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0101111100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1737|picorv32_core/reg15_b35  (
    .a({\picorv32_core/n667_lutinv ,_al_u1735_o}),
    .b({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdcycleh }),
    .c({_al_u1313_o,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1736_o,\picorv32_core/count_cycle [35]}),
    .e({\picorv32_core/pcpi_rs1$3$ ,\picorv32_core/count_instr [3]}),
    .mi({open_n9108,\picorv32_core/n459 [35]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1737_o,_al_u1736_o}),
    .q({open_n9123,\picorv32_core/count_cycle [35]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0010101000101010),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u1738|_al_u1860  (
    .a({open_n9124,_al_u1859_o}),
    .b({\picorv32_core/n666_lutinv ,\picorv32_core/n666_lutinv }),
    .c({\picorv32_core/n543 [3],\picorv32_core/n543 [14]}),
    .d({_al_u1737_o,open_n9127}),
    .f({_al_u1738_o,_al_u1860_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)"),
    //.LUT1("(C*B*A)"),
    .INIT_LUT0(16'b1100110010101010),
    .INIT_LUT1(16'b1000000010000000),
    .MODE("LOGIC"))
    \_al_u1740|_al_u1521  (
    .a({mem_rdata[29],memory_out[29]}),
    .b({\picorv32_core/n734_lutinv ,uart_do[29]}),
    .c({\picorv32_core/latched_is_lu ,open_n9146}),
    .d({open_n9149,uart_sel_lutinv_placeOpt_1}),
    .f({\picorv32_core/sel27_b29/B2 ,mem_rdata[29]}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("(~B*~D*~(0*~(A*~C)))"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("(~B*~D*~(1*~(A*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1741|picorv32_core/reg13_b29  (
    .a({_al_u1661_o,_al_u1745_o}),
    .b({\picorv32_core/sel27_b29/B2 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .c({_al_u1658_o,_al_u1741_o}),
    .clk(clk_pad),
    .d({\picorv32_core/sel27_b16/B1 ,\picorv32_core/n580 }),
    .e({\picorv32_core/latched_is_lb ,resetn_placeOpt_13}),
    .f({_al_u1741_o,open_n9184}),
    .q({open_n9188,\picorv32_core/reg_out [29]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~C*~(0*A)*~(~D*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~C*~(1*A)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000111100000011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000010100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1745|picorv32_core/reg15_b61  (
    .a({\picorv32_core/n666_lutinv ,_al_u1743_o}),
    .b({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdcycleh }),
    .c({\picorv32_core/sel43_b29/B2 ,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1744_o,\picorv32_core/count_cycle [61]}),
    .e({\picorv32_core/n543 [29],\picorv32_core/count_instr [29]}),
    .mi({open_n9191,\picorv32_core/n459 [61]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1745_o,_al_u1744_o}),
    .q({open_n9206,\picorv32_core/count_cycle [61]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    //.LUT1("(D*C*B)"),
    .INIT_LUT0(16'b1010101011001100),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1747|_al_u1523  (
    .a({open_n9207,uart_do[28]}),
    .b({mem_rdata[28],memory_out[28]}),
    .c({\picorv32_core/n734_lutinv ,open_n9208}),
    .d({\picorv32_core/latched_is_lu ,uart_sel_lutinv_placeOpt_1}),
    .f({\picorv32_core/sel27_b28/B2 ,mem_rdata[28]}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("(~B*~A*~(0*~(C*~D)))"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("(~B*~A*~(1*~(C*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1748|picorv32_core/reg13_b28  (
    .a({\picorv32_core/sel27_b16/B1 ,_al_u1752_o}),
    .b({\picorv32_core/sel27_b28/B2 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .c({_al_u1661_o,_al_u1748_o}),
    .clk(clk_pad),
    .d({_al_u1658_o,\picorv32_core/n580 }),
    .e({\picorv32_core/latched_is_lb ,resetn_placeOpt_13}),
    .f({_al_u1748_o,open_n9245}),
    .q({open_n9249,\picorv32_core/reg_out [28]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~C*~(0*A)*~(~D*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~C*~(1*A)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000111100000011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000010100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1752|picorv32_core/reg15_b28  (
    .a({\picorv32_core/n666_lutinv ,_al_u1750_o}),
    .b({\picorv32_core/n664_lutinv_placeOpt_1 ,\picorv32_core/instr_rdcycle }),
    .c({\picorv32_core/sel43_b28/B2 ,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1751_o,\picorv32_core/count_cycle [28]}),
    .e({\picorv32_core/n543 [28],\picorv32_core/count_instr [60]}),
    .mi({open_n9252,\picorv32_core/n459 [28]}),
    .sr(resetn_placeOpt_8),
    .f({_al_u1752_o,_al_u1751_o}),
    .q({open_n9267,\picorv32_core/count_cycle [28]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~B*~(0*~(C*~D)))"),
    //.LUTF1("(B*D*A)"),
    //.LUTG0("(~A*~B*~(1*~(C*~D)))"),
    //.LUTG1("(B*D*A)"),
    .INIT_LUTF0(16'b0001000100010001),
    .INIT_LUTF1(16'b1000100000000000),
    .INIT_LUTG0(16'b0000000000010000),
    .INIT_LUTG1(16'b1000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1754|_al_u1755  (
    .a({mem_rdata[27],\picorv32_core/sel27_b27/B2 }),
    .b({\picorv32_core/latched_is_lu ,\picorv32_core/sel27_b16/B1 }),
    .c({open_n9268,_al_u1661_o}),
    .d({\picorv32_core/n734_lutinv ,_al_u1658_o}),
    .e({open_n9271,\picorv32_core/latched_is_lb }),
    .f({\picorv32_core/sel27_b27/B2 ,_al_u1755_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1758|picorv32_core/reg15_b59  (
    .a({_al_u1757_o,_al_u1756_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycleh }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [59]}),
    .e({\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/count_instr [27]}),
    .mi({open_n9294,\picorv32_core/n459 [59]}),
    .sr(resetn_placeOpt_9),
    .f({_al_u1758_o,_al_u1757_o}),
    .q({open_n9309,\picorv32_core/count_cycle [59]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C*D))"),
    //.LUT1("(D*~(A*C))"),
    .INIT_LUT0(16'b0000101010101010),
    .INIT_LUT1(16'b0101111100000000),
    .MODE("LOGIC"))
    \_al_u1759|_al_u1853  (
    .a({\picorv32_core/n543 [27],_al_u1852_o}),
    .c({\picorv32_core/n666_lutinv ,\picorv32_core/n543 [15]}),
    .d({_al_u1758_o,\picorv32_core/n666_lutinv }),
    .f({_al_u1759_o,_al_u1853_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1010000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1761|_al_u1812  (
    .a({open_n9332,\picorv32_core/pcpi_rs1$1$ }),
    .b({\picorv32_core/n734_lutinv ,open_n9333}),
    .c({\picorv32_core/latched_is_lu ,\picorv32_core/pcpi_rs1$0$ }),
    .d({mem_rdata[26],mem_rdata[26]}),
    .f({\picorv32_core/sel27_b26/B2 ,_al_u1812_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B*~(0*~(C*~D)))"),
    //.LUT1("(~A*~B*~(1*~(C*~D)))"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0000000000010000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1762 (
    .a({\picorv32_core/sel27_b26/B2 ,\picorv32_core/sel27_b26/B2 }),
    .b({\picorv32_core/sel27_b16/B1 ,\picorv32_core/sel27_b16/B1 }),
    .c({_al_u1661_o,_al_u1661_o}),
    .d({_al_u1658_o,_al_u1658_o}),
    .mi({open_n9366,\picorv32_core/latched_is_lb }),
    .fx({open_n9371,_al_u1762_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*C*A)*~(~D*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*C*A)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1111111100110011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0101111100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1765|picorv32_core/reg15_b26  (
    .a({\picorv32_core/n667_lutinv ,_al_u1763_o}),
    .b({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdcycle }),
    .c({_al_u1313_o,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1764_o,\picorv32_core/count_cycle [26]}),
    .e({\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/count_instr [58]}),
    .mi({open_n9376,\picorv32_core/n459 [26]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1765_o,_al_u1764_o}),
    .q({open_n9391,\picorv32_core/count_cycle [26]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~D*~B*C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    //.LUTF1("~B*~A*~C*D+B*~A*~C*D+~B*A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG0("~A*~D*~B*C+A*~D*~B*C+~A*~D*B*C+A*~D*B*C"),
    //.LUTG1("~B*~A*~C*D+B*~A*~C*D+~B*~A*C*D+B*~A*C*D"),
    .INIT_LUTF0(16'b1111000011110000),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0101010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1766|_al_u1846  (
    .a({\picorv32_core/n666_lutinv ,open_n9392}),
    .c({open_n9395,_al_u1845_o}),
    .d({_al_u1765_o,\picorv32_core/n666_lutinv }),
    .e({\picorv32_core/n543 [26],\picorv32_core/n543 [16]}),
    .f({_al_u1766_o,_al_u1846_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("(~B*~C*~(0*~(A*~D)))"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("(~B*~C*~(1*~(A*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000001100000011),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1769|picorv32_core/reg13_b25  (
    .a({_al_u1661_o,_al_u1773_o}),
    .b({\picorv32_core/sel27_b25/B2 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .c({\picorv32_core/sel27_b16/B1 ,_al_u1769_o}),
    .clk(clk_pad),
    .d({_al_u1658_o,\picorv32_core/n580 }),
    .e({\picorv32_core/latched_is_lb ,resetn_placeOpt_13}),
    .f({_al_u1769_o,open_n9434}),
    .q({open_n9438,\picorv32_core/reg_out [25]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1772|picorv32_core/reg15_b57  (
    .a({_al_u1771_o,_al_u1770_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycleh }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [57]}),
    .e({\picorv32_core/pcpi_rs1$25$ ,\picorv32_core/count_instr [25]}),
    .mi({open_n9441,\picorv32_core/n459 [57]}),
    .sr(resetn_placeOpt_4),
    .f({_al_u1772_o,_al_u1771_o}),
    .q({open_n9456,\picorv32_core/count_cycle [57]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~D*~B*C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    //.LUTF1("~B*~D*~C*A+B*~D*~C*A+~B*D*~C*A+B*D*~C*A+~B*~D*C*A+B*~D*C*A+~B*D*C*A+B*D*C*A"),
    //.LUTG0("~A*~D*~B*C+A*~D*~B*C+~A*~D*B*C+A*~D*B*C"),
    //.LUTG1("~B*~D*~C*A+B*~D*~C*A+~B*~D*C*A+B*~D*C*A"),
    .INIT_LUTF0(16'b1111000011110000),
    .INIT_LUTF1(16'b1010101010101010),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1773|_al_u1839  (
    .a({_al_u1772_o,open_n9457}),
    .c({open_n9460,_al_u1838_o}),
    .d({\picorv32_core/n666_lutinv ,\picorv32_core/n666_lutinv }),
    .e({\picorv32_core/n543 [25],\picorv32_core/n543 [17]}),
    .f({_al_u1773_o,_al_u1839_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*C*~D+A*B*C*~D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("(D*C*A)"),
    //.LUTG0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("(D*C*A)"),
    .INIT_LUTF0(16'b1010000010100000),
    .INIT_LUTF1(16'b1010000000000000),
    .INIT_LUTG0(16'b1111010111110101),
    .INIT_LUTG1(16'b1010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1775|_al_u1503  (
    .a({mem_rdata[24],uart_sel_lutinv_placeOpt_3}),
    .c({\picorv32_core/n734_lutinv ,uart_do[24]}),
    .d({\picorv32_core/latched_is_lu ,open_n9487}),
    .e({open_n9488,memory_out[24]}),
    .f({\picorv32_core/sel27_b24/B2 ,mem_rdata[24]}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("(~B*~D*~(0*~(A*~C)))"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("(~B*~D*~(1*~(A*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1776|picorv32_core/reg13_b24  (
    .a({_al_u1661_o,_al_u1780_o}),
    .b({\picorv32_core/sel27_b24/B2 ,\picorv32_core/n669_lutinv }),
    .c({_al_u1658_o,_al_u1776_o}),
    .clk(clk_pad),
    .d({\picorv32_core/sel27_b16/B1 ,\picorv32_core/n580 }),
    .e({\picorv32_core/latched_is_lb ,resetn_placeOpt_10}),
    .f({_al_u1776_o,open_n9525}),
    .q({open_n9529,\picorv32_core/reg_out [24]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*C*A)*~(~D*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*C*A)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1111111100110011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0101111100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1779|picorv32_core/reg15_b56  (
    .a({\picorv32_core/n667_lutinv ,_al_u1777_o}),
    .b({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdcycleh }),
    .c({_al_u1313_o,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1778_o,\picorv32_core/count_cycle [56]}),
    .e({\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/count_instr [24]}),
    .mi({open_n9532,\picorv32_core/n459 [56]}),
    .sr(resetn_placeOpt_9),
    .f({_al_u1779_o,_al_u1778_o}),
    .q({open_n9547,\picorv32_core/count_cycle [56]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(C*~(A*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0111000001110000),
    .MODE("LOGIC"))
    \_al_u1780|_al_u1832  (
    .a({\picorv32_core/n543 [24],open_n9548}),
    .b({\picorv32_core/n666_lutinv ,\picorv32_core/n666_lutinv }),
    .c({_al_u1779_o,\picorv32_core/n543 [18]}),
    .d({open_n9551,_al_u1831_o}),
    .f({_al_u1780_o,_al_u1832_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*A)"),
    //.LUT1("(D*B*C)"),
    .INIT_LUT0(16'b1000000010000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1782|_al_u1768  (
    .a({open_n9570,mem_rdata[25]}),
    .b({\picorv32_core/n734_lutinv ,\picorv32_core/n734_lutinv }),
    .c({mem_rdata[23],\picorv32_core/latched_is_lu }),
    .d({\picorv32_core/latched_is_lu ,open_n9573}),
    .f({\picorv32_core/sel27_b23/B2 ,\picorv32_core/sel27_b25/B2 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B*~(0*~(C*~D)))"),
    //.LUT1("(~B*~C*~(1*~(D*~A)))"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0000000100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1783 (
    .a({_al_u1658_o,\picorv32_core/sel27_b23/B2 }),
    .b({\picorv32_core/sel27_b23/B2 ,\picorv32_core/sel27_b16/B1 }),
    .c({\picorv32_core/sel27_b16/B1 ,_al_u1661_o}),
    .d({_al_u1661_o,_al_u1658_o}),
    .mi({open_n9604,\picorv32_core/latched_is_lb }),
    .fx({open_n9609,_al_u1783_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1786|picorv32_core/reg15_b55  (
    .a({_al_u1785_o,_al_u1784_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycleh }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [55]}),
    .e({\picorv32_core/pcpi_rs1$23$ ,\picorv32_core/count_instr [23]}),
    .mi({open_n9614,\picorv32_core/n459 [55]}),
    .sr(resetn_placeOpt_9),
    .f({_al_u1786_o,_al_u1785_o}),
    .q({open_n9629,\picorv32_core/count_cycle [55]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*D))"),
    //.LUT1("(C*~(A*D))"),
    .INIT_LUT0(16'b0101000011110000),
    .INIT_LUT1(16'b0101000011110000),
    .MODE("LOGIC"))
    \_al_u1787|_al_u1825  (
    .a({\picorv32_core/n543 [23],\picorv32_core/n543 [19]}),
    .c({_al_u1786_o,_al_u1824_o}),
    .d({\picorv32_core/n666_lutinv ,\picorv32_core/n666_lutinv }),
    .f({_al_u1787_o,_al_u1825_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~B*~(0*~(C*~D)))"),
    //.LUTF1("0"),
    //.LUTG0("(~A*~B*~(1*~(C*~D)))"),
    //.LUTG1("~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0001000100010001),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000010000),
    .INIT_LUTG1(16'b1100110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1789|_al_u1790  (
    .a({open_n9652,\picorv32_core/sel27_b22/B2 }),
    .b({\picorv32_core/latched_is_lu ,\picorv32_core/sel27_b16/B1 }),
    .c({open_n9653,_al_u1661_o}),
    .d({mem_rdata[22],_al_u1658_o}),
    .e({\picorv32_core/n734_lutinv ,\picorv32_core/latched_is_lb }),
    .f({\picorv32_core/sel27_b22/B2 ,_al_u1790_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*C*A)*~(~D*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*C*A)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1111111100110011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0101111100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1793|picorv32_core/reg15_b54  (
    .a({\picorv32_core/n667_lutinv ,_al_u1791_o}),
    .b({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdcycleh }),
    .c({_al_u1313_o,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1792_o,\picorv32_core/count_cycle [54]}),
    .e({\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/count_instr [22]}),
    .mi({open_n9678,\picorv32_core/n459 [54]}),
    .sr(resetn_placeOpt_4),
    .f({_al_u1793_o,_al_u1792_o}),
    .q({open_n9693,\picorv32_core/count_cycle [54]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D+A*~B*~C*D+A*B*~C*D"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*~C*D+A*B*~C*D"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b1010101010101010),
    .INIT_LUTG0(16'b0000101000001010),
    .INIT_LUTG1(16'b0000101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1794|_al_u1818  (
    .a({_al_u1793_o,_al_u1817_o}),
    .c({\picorv32_core/n543 [22],\picorv32_core/n543 [2]}),
    .e({\picorv32_core/n666_lutinv ,\picorv32_core/n666_lutinv }),
    .f({_al_u1794_o,_al_u1818_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTF1("(D*B*A)"),
    //.LUTG0("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("(D*B*A)"),
    .INIT_LUTF0(16'b0000000011001100),
    .INIT_LUTF1(16'b1000100000000000),
    .INIT_LUTG0(16'b1111111111001100),
    .INIT_LUTG1(16'b1000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1796|_al_u1509  (
    .a({mem_rdata[21],open_n9720}),
    .b({\picorv32_core/n734_lutinv ,memory_out[21]}),
    .d({\picorv32_core/latched_is_lu ,uart_sel_lutinv_placeOpt_1}),
    .e({open_n9725,uart_do[21]}),
    .f({\picorv32_core/sel27_b21/B2 ,mem_rdata[21]}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("(~B*~A*~(0*~(D*~C)))"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("(~B*~A*~(1*~(D*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1797|picorv32_core/reg13_b21  (
    .a({\picorv32_core/sel27_b16/B1 ,_al_u1801_o}),
    .b({\picorv32_core/sel27_b21/B2 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .c({_al_u1658_o,_al_u1797_o}),
    .clk(clk_pad),
    .d({_al_u1661_o,\picorv32_core/n580 }),
    .e({\picorv32_core/latched_is_lb ,resetn_placeOpt_13}),
    .f({_al_u1797_o,open_n9762}),
    .q({open_n9766,\picorv32_core/reg_out [21]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0111111101111111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0111111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1800|picorv32_core/reg15_b53  (
    .a({\picorv32_core/n667_lutinv ,_al_u1798_o}),
    .b({\picorv32_core/pcpi_rs1$21$ ,\picorv32_core/instr_rdcycleh }),
    .c({_al_u1313_o,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1799_o,\picorv32_core/count_cycle [53]}),
    .e({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/count_instr [21]}),
    .mi({open_n9769,\picorv32_core/n459 [53]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1800_o,_al_u1799_o}),
    .q({open_n9784,\picorv32_core/count_cycle [53]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~D*~B*C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    //.LUTF1("~A*~D*~B*C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    //.LUTG0("~A*~D*~B*C+A*~D*~B*C+~A*~D*B*C+A*~D*B*C"),
    //.LUTG1("~A*~D*~B*C+A*~D*~B*C+~A*~D*B*C+A*~D*B*C"),
    .INIT_LUTF0(16'b1111000011110000),
    .INIT_LUTF1(16'b1111000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1801|_al_u1808  (
    .c({_al_u1800_o,_al_u1807_o}),
    .d({\picorv32_core/n666_lutinv ,\picorv32_core/n666_lutinv }),
    .e(\picorv32_core/n543 [21:20]),
    .f({_al_u1801_o,_al_u1808_o}));
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTF1("0"),
    //.LUTG0("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTG1("~C*A*B*~D+C*A*B*~D+~C*A*B*D+C*A*B*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010011000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1110111011001111),
    .INIT_LUTG1(16'b1000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1803|picorv32_core/reg5_b4  (
    .a({\picorv32_core/n734_lutinv ,_al_u1089_o}),
    .b({\picorv32_core/latched_is_lu ,mem_rdata[20]}),
    .c({open_n9811,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({open_n9812,\picorv32_core/mem_la_read }),
    .e({mem_rdata[20],\picorv32_core/mem_16bit_buffer [4]}),
    .f({\picorv32_core/sel27_b20/B2 ,open_n9828}),
    .q({open_n9832,\picorv32_core/mem_16bit_buffer [4]}));  // ../src/picorv32.v(605)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("(~C*~A*~(0*~(B*~D)))"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("(~C*~A*~(1*~(B*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000010100000101),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1804|picorv32_core/reg13_b20  (
    .a({\picorv32_core/sel27_b16/B1 ,_al_u1808_o}),
    .b({_al_u1661_o,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .c({\picorv32_core/sel27_b20/B2 ,_al_u1804_o}),
    .clk(clk_pad),
    .d({_al_u1658_o,\picorv32_core/n580 }),
    .e({\picorv32_core/latched_is_lb ,resetn_placeOpt_13}),
    .f({_al_u1804_o,open_n9849}),
    .q({open_n9853,\picorv32_core/reg_out [20]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1807|picorv32_core/reg15_b20  (
    .a({_al_u1806_o,_al_u1805_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycle }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [20]}),
    .e({\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/count_instr [52]}),
    .mi({open_n9856,\picorv32_core/n459 [20]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1807_o,_al_u1806_o}),
    .q({open_n9871,\picorv32_core/count_cycle [20]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~((B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D))*~(C)+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*~(C)+~(A)*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C+A*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)*C)"),
    //.LUTF1("A*B*~C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("(A*~((B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D))*~(C)+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*~(C)+~(A)*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C+A*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)*C)"),
    //.LUTG1("A*B*~C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000101011001010),
    .INIT_LUTF1(16'b1011101110001000),
    .INIT_LUTG0(16'b1111101011001010),
    .INIT_LUTG1(16'b1011101110001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1810|_al_u1269  (
    .a({uart_do[2],\picorv32_core/mem_rdata_q [2]}),
    .b({uart_sel_lutinv_placeOpt_2,memory_out[2]}),
    .c({open_n9872,\picorv32_core/mem_xfer_placeOpt_4 }),
    .d({memory_out[2],uart_sel_lutinv_placeOpt_2}),
    .e({open_n9875,uart_do[2]}),
    .f({mem_rdata[2],\picorv32_core/mem_rdata_latched_noshuffle [2]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D)"),
    //.LUT1("(~(A*C)*~(~B*D))"),
    .INIT_LUT0(16'b1111000010101010),
    .INIT_LUT1(16'b0100110001011111),
    .MODE("LOGIC"))
    \_al_u1811|_al_u1515  (
    .a({_al_u1660_o,memory_out[18]}),
    .b({_al_u1136_o,open_n9896}),
    .c({mem_rdata[18],uart_do[18]}),
    .d({mem_rdata[2],uart_sel_lutinv_placeOpt_1}),
    .f({_al_u1811_o,mem_rdata[18]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(D*~(0*~(~B*~(A*C))))"),
    //.LUTG0("(~1*~B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(D*~(1*~(~B*~(A*C))))"),
    .INIT_LUTF0(16'b0010001100100000),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0001001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1814|_al_u1883  (
    .a({\picorv32_core/n40 [1],mem_rdata[26]}),
    .b({_al_u1812_o,\picorv32_core/latched_is_lb }),
    .c({mem_rdata[10],_al_u1663_o}),
    .d({_al_u1811_o,mem_rdata[10]}),
    .e({_al_u1657_o,\picorv32_core/mem_wordsize [1]}),
    .f({_al_u1814_o,_al_u1883_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*C*A)*~(~D*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*C*A)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1111111100110011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0101111100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1817|picorv32_core/reg15_b34  (
    .a({\picorv32_core/n667_lutinv ,_al_u1815_o}),
    .b({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdcycleh }),
    .c({_al_u1313_o,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1816_o,\picorv32_core/count_cycle [34]}),
    .e({\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/count_instr [2]}),
    .mi({open_n9941,\picorv32_core/n459 [34]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1817_o,_al_u1816_o}),
    .q({open_n9956,\picorv32_core/count_cycle [34]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~C*~(0*~(B*~D)))"),
    //.LUTF1("0"),
    //.LUTG0("(~A*~C*~(1*~(B*~D)))"),
    //.LUTG1("~B*C*A*~D+B*C*A*~D+~B*C*A*D+B*C*A*D"),
    .INIT_LUTF0(16'b0000010100000101),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000100),
    .INIT_LUTG1(16'b1010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1820|_al_u1821  (
    .a({\picorv32_core/latched_is_lu ,\picorv32_core/sel27_b19/B2 }),
    .b({open_n9957,_al_u1661_o}),
    .c({\picorv32_core/n734_lutinv ,\picorv32_core/sel27_b16/B1 }),
    .d({open_n9960,_al_u1658_o}),
    .e({mem_rdata[19],\picorv32_core/latched_is_lb }),
    .f({\picorv32_core/sel27_b19/B2 ,_al_u1821_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1824|picorv32_core/reg15_b19  (
    .a({_al_u1823_o,_al_u1822_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycle }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [19]}),
    .e({\picorv32_core/pcpi_rs1$19$ ,\picorv32_core/count_instr [51]}),
    .mi({open_n9983,\picorv32_core/n459 [19]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1824_o,_al_u1823_o}),
    .q({open_n9998,\picorv32_core/count_cycle [19]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("(~B*~D*~(0*~(A*~C)))"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("(~B*~D*~(1*~(A*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1828|picorv32_core/reg13_b18  (
    .a({_al_u1661_o,_al_u1832_o}),
    .b({\picorv32_core/sel27_b18/B2 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .c({_al_u1658_o,_al_u1828_o}),
    .clk(clk_pad),
    .d({\picorv32_core/sel27_b16/B1 ,\picorv32_core/n580 }),
    .e({\picorv32_core/latched_is_lb ,resetn_placeOpt_12}),
    .f({_al_u1828_o,open_n10015}),
    .q({open_n10019,\picorv32_core/reg_out [18]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1831|picorv32_core/reg15_b18  (
    .a({_al_u1830_o,_al_u1829_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycle }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [18]}),
    .e({\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/count_instr [50]}),
    .mi({open_n10022,\picorv32_core/n459 [18]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1831_o,_al_u1830_o}),
    .q({open_n10037,\picorv32_core/count_cycle [18]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D)"),
    //.LUTF1("0"),
    //.LUTG0("(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D)"),
    //.LUTG1("A*D*~C*~B+A*D*C*~B+A*D*~C*B+A*D*C*B"),
    .INIT_LUTF0(16'b1111000010101010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010101010),
    .INIT_LUTG1(16'b1010101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1834|_al_u1528  (
    .a({mem_rdata[17],memory_out[17]}),
    .c({open_n10040,uart_do[17]}),
    .d({\picorv32_core/n734_lutinv ,uart_sel_lutinv_placeOpt_1}),
    .e({\picorv32_core/latched_is_lu ,open_n10043}),
    .f({\picorv32_core/sel27_b17/B2 ,mem_rdata[17]}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("(~B*~D*~(0*~(A*~C)))"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("(~B*~D*~(1*~(A*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1835|picorv32_core/reg13_b17  (
    .a({_al_u1661_o,_al_u1839_o}),
    .b({\picorv32_core/sel27_b17/B2 ,\picorv32_core/n669_lutinv }),
    .c({_al_u1658_o,_al_u1835_o}),
    .clk(clk_pad),
    .d({\picorv32_core/sel27_b16/B1 ,\picorv32_core/n580 }),
    .e({\picorv32_core/latched_is_lb ,resetn_placeOpt_10}),
    .f({_al_u1835_o,open_n10080}),
    .q({open_n10084,\picorv32_core/reg_out [17]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1838|picorv32_core/reg15_b49  (
    .a({_al_u1837_o,_al_u1836_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycleh }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [49]}),
    .e({\picorv32_core/pcpi_rs1$17$ ,\picorv32_core/count_instr [17]}),
    .mi({open_n10087,\picorv32_core/n459 [49]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1838_o,_al_u1837_o}),
    .q({open_n10102,\picorv32_core/count_cycle [49]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(605)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTF1("(A*B*C)"),
    //.LUTG0("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUTG1("(A*B*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010011000000),
    .INIT_LUTF1(16'b1000000010000000),
    .INIT_LUTG0(16'b1110111011001111),
    .INIT_LUTG1(16'b1000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1841|picorv32_core/reg5_b0  (
    .a({\picorv32_core/latched_is_lu ,_al_u1089_o}),
    .b({\picorv32_core/n734_lutinv ,mem_rdata[16]}),
    .c({mem_rdata[16],\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({open_n10103,\picorv32_core/mem_la_read }),
    .e({open_n10104,\picorv32_core/mem_16bit_buffer [0]}),
    .f({\picorv32_core/sel27_b16/B2 ,open_n10120}),
    .q({open_n10124,\picorv32_core/mem_16bit_buffer [0]}));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~C*~(0*~(B*~D)))"),
    //.LUT1("(~A*~C*~(1*~(B*~D)))"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1842 (
    .a({\picorv32_core/sel27_b16/B2 ,\picorv32_core/sel27_b16/B2 }),
    .b({_al_u1661_o,_al_u1661_o}),
    .c({\picorv32_core/sel27_b16/B1 ,\picorv32_core/sel27_b16/B1 }),
    .d({_al_u1658_o,_al_u1658_o}),
    .mi({open_n10137,\picorv32_core/latched_is_lb }),
    .fx({open_n10142,_al_u1842_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1845|picorv32_core/reg15_b16  (
    .a({_al_u1844_o,_al_u1843_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycle }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [16]}),
    .e({\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/count_instr [48]}),
    .mi({open_n10147,\picorv32_core/n459 [16]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1845_o,_al_u1844_o}),
    .q({open_n10162,\picorv32_core/count_cycle [16]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(A*C*D)"),
    //.LUT1("(~C*~(A*B))"),
    .INIT_LUT0(16'b1010000000000000),
    .INIT_LUT1(16'b0000011100000111),
    .MODE("LOGIC"))
    \_al_u1848|_al_u1715  (
    .a({_al_u1713_o,\picorv32_core/latched_is_lu }),
    .b({mem_rdata[31],open_n10163}),
    .c({_al_u1712_o,\picorv32_core/n734_lutinv }),
    .d({open_n10166,mem_rdata[31]}),
    .f({_al_u1848_o,\picorv32_core/sel27_b31/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*~D*~A+~C*B*~D*~A+~C*~B*~D*A+~C*B*~D*A"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("~C*~B*~D*~A+C*~B*~D*~A+~C*B*~D*~A+~C*~B*~D*A+C*~B*~D*A+~C*B*~D*A"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1011111110111111),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1000110010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1849|_al_u1870  (
    .a({_al_u1658_o,open_n10185}),
    .b({\picorv32_core/latched_is_lb ,_al_u1658_o}),
    .c({_al_u1661_o,\picorv32_core/latched_is_lb }),
    .d({open_n10188,_al_u1869_o}),
    .e({_al_u1848_o,_al_u1661_o}),
    .f({_al_u1849_o,_al_u1870_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1852|picorv32_core/reg15_b47  (
    .a({_al_u1851_o,_al_u1850_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycleh }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [47]}),
    .e({\picorv32_core/pcpi_rs1$15$ ,\picorv32_core/count_instr [15]}),
    .mi({open_n10211,\picorv32_core/n459 [47]}),
    .sr(resetn_placeOpt_4),
    .f({_al_u1852_o,_al_u1851_o}),
    .q({open_n10226,\picorv32_core/count_cycle [47]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("~B*~C*~A*~D+B*~C*~A*~D+~B*~C*A*~D+B*~C*A*~D+~B*C*A*~D+B*C*A*~D"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("~B*~C*~A*~D+B*~C*~A*~D+~B*~C*A*~D+B*~C*A*~D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000010101111),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1856|picorv32_core/reg13_b14  (
    .a({_al_u1661_o,_al_u1860_o}),
    .b({open_n10227,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .c({\picorv32_core/latched_is_lb ,_al_u1856_o}),
    .clk(clk_pad),
    .d({_al_u1855_o,\picorv32_core/n580 }),
    .e({_al_u1658_o,resetn_placeOpt_12}),
    .f({_al_u1856_o,open_n10244}),
    .q({open_n10248,\picorv32_core/reg_out [14]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*D*B)*~(~A*C))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1859|picorv32_core/reg15_b14  (
    .a({_al_u1858_o,_al_u1857_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycle }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [14]}),
    .e({\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/count_instr [46]}),
    .mi({open_n10251,\picorv32_core/n459 [14]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1859_o,_al_u1858_o}),
    .q({open_n10266,\picorv32_core/count_cycle [14]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("~C*~B*~A*~D+~C*~B*A*~D+~C*~B*~A*D+~C*~B*A*D"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("~C*~B*~A*~D+~C*B*~A*~D+~C*~B*A*~D+~C*B*A*~D+~C*~B*~A*D+~C*~B*A*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000001100000011),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1863|picorv32_core/reg13_b13  (
    .a({open_n10267,_al_u1867_o}),
    .b({\picorv32_core/latched_is_lb ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .c({_al_u1862_o,_al_u1863_o}),
    .clk(clk_pad),
    .d({_al_u1658_o,\picorv32_core/n580 }),
    .e({_al_u1661_o,resetn_placeOpt_12}),
    .f({_al_u1863_o,open_n10284}),
    .q({open_n10288,\picorv32_core/reg_out [13]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*C*A)*~(~D*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*C*A)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1111111100110011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0101111100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1866|picorv32_core/reg15_b13  (
    .a({\picorv32_core/n667_lutinv ,_al_u1864_o}),
    .b({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdcycle }),
    .c({_al_u1313_o,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1865_o,\picorv32_core/count_cycle [13]}),
    .e({\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/count_instr [45]}),
    .mi({open_n10291,\picorv32_core/n459 [13]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1866_o,_al_u1865_o}),
    .q({open_n10306,\picorv32_core/count_cycle [13]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~1*~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1869 (
    .a({_al_u1663_o,\picorv32_core/latched_is_lb }),
    .b({\picorv32_core/latched_is_lb ,_al_u1663_o}),
    .c({mem_rdata[12],mem_rdata[12]}),
    .d({mem_rdata[28],mem_rdata[28]}),
    .mi({open_n10319,\picorv32_core/mem_wordsize [1]}),
    .fx({open_n10324,_al_u1869_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*C*A)*~(~D*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*C*A)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1111111100110011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0101111100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1873|picorv32_core/reg15_b44  (
    .a({\picorv32_core/n667_lutinv ,_al_u1871_o}),
    .b({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdcycleh }),
    .c({_al_u1313_o,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1872_o,\picorv32_core/count_cycle [44]}),
    .e({\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/count_instr [12]}),
    .mi({open_n10329,\picorv32_core/n459 [44]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1873_o,_al_u1872_o}),
    .q({open_n10344,\picorv32_core/count_cycle [44]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("(~1*~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUT0(16'b0010001100100000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1876 (
    .a({_al_u1663_o,mem_rdata[27]}),
    .b({\picorv32_core/latched_is_lb ,\picorv32_core/latched_is_lb }),
    .c({mem_rdata[11],_al_u1663_o}),
    .d({mem_rdata[27],mem_rdata[11]}),
    .mi({open_n10357,\picorv32_core/mem_wordsize [1]}),
    .fx({open_n10362,_al_u1876_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1880|picorv32_core/reg15_b43  (
    .a({_al_u1879_o,_al_u1878_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/instr_rdcycleh }),
    .c({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1313_o,\picorv32_core/count_cycle [43]}),
    .e({\picorv32_core/pcpi_rs1$11$ ,\picorv32_core/count_instr [11]}),
    .mi({open_n10367,\picorv32_core/n459 [43]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1880_o,_al_u1879_o}),
    .q({open_n10382,\picorv32_core/count_cycle [43]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("~A*~B*C*~D+~A*B*C*~D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1884|picorv32_core/reg13_b10  (
    .a({_al_u1883_o,_al_u1888_o}),
    .b({open_n10383,\picorv32_core/n669_lutinv }),
    .c({_al_u1661_o,_al_u1884_o}),
    .clk(clk_pad),
    .d({_al_u1658_o,\picorv32_core/n580 }),
    .e({\picorv32_core/latched_is_lb ,resetn_placeOpt_10}),
    .f({_al_u1884_o,open_n10400}),
    .q({open_n10404,\picorv32_core/reg_out [10]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*C*A)*~(~D*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*C*A)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1111111100110011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0101111100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1887|picorv32_core/reg15_b10  (
    .a({\picorv32_core/n667_lutinv ,_al_u1885_o}),
    .b({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdcycle }),
    .c({_al_u1313_o,\picorv32_core/instr_rdinstrh }),
    .clk(clk_pad),
    .d({_al_u1886_o,\picorv32_core/count_cycle [10]}),
    .e({\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/count_instr [42]}),
    .mi({open_n10407,\picorv32_core/n459 [10]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1887_o,_al_u1886_o}),
    .q({open_n10422,\picorv32_core/count_cycle [10]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*(C*~(D)*~(0)+C*D*~(0)+~(C)*D*0+C*D*0))"),
    //.LUT1("(B*A*(C*~(D)*~(1)+C*D*~(1)+~(C)*D*1+C*D*1))"),
    .INIT_LUT0(16'b1000000010000000),
    .INIT_LUT1(16'b1000100000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1890 (
    .a({_al_u1657_o,_al_u1657_o}),
    .b({\picorv32_core/pcpi_rs1$0$ ,\picorv32_core/pcpi_rs1$0$ }),
    .c({mem_rdata[9],mem_rdata[9]}),
    .d({mem_rdata[25],mem_rdata[25]}),
    .mi({open_n10435,\picorv32_core/pcpi_rs1$1$ }),
    .fx({open_n10440,_al_u1890_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(A*~(B*~C*D)))"),
    //.LUTF1("(~C*~(~B*A)*~(0*D))"),
    //.LUTG0("(1*~(A*~(B*~C*D)))"),
    //.LUTG1("(~C*~(~B*A)*~(1*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000110100001101),
    .INIT_LUTG0(16'b0101110101010101),
    .INIT_LUTG1(16'b0000000000001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1891|picorv32_core/reg13_b1  (
    .a({mem_rdata[1],_al_u1895_o}),
    .b({_al_u1136_o,\picorv32_core/n669_lutinv }),
    .c({_al_u1890_o,_al_u1891_o}),
    .clk(clk_pad),
    .d({mem_rdata[17],\picorv32_core/n580 }),
    .e({_al_u1660_o,resetn_placeOpt_10}),
    .f({_al_u1891_o,open_n10459}),
    .q({open_n10463,\picorv32_core/reg_out [1]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~(0*C*A)*~(~D*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~(1*C*A)*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1111111100110011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0101111100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1894|picorv32_core/reg19_b33  (
    .a({\picorv32_core/n667_lutinv ,_al_u1892_o}),
    .b({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdcycle }),
    .c({_al_u1313_o,\picorv32_core/instr_rdinstrh }),
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({_al_u1893_o,\picorv32_core/count_cycle [1]}),
    .e({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/count_instr [33]}),
    .mi({open_n10465,\picorv32_core/n503 [33]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1894_o,_al_u1893_o}),
    .q({open_n10480,\picorv32_core/count_instr [33]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(B*D)*~(~A*C))"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"))
    \_al_u1898|_al_u1897  (
    .a({_al_u1136_o,open_n10481}),
    .b({_al_u1660_o,memory_out[0]}),
    .c({mem_rdata[0],uart_do[0]}),
    .d({mem_rdata[16],uart_sel_lutinv}),
    .f({_al_u1898_o,mem_rdata[0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(0*~(~C*~(A*B))))"),
    //.LUT1("(D*~(1*~(~C*~(A*B))))"),
    .INIT_LUT0(16'b1111111100000000),
    .INIT_LUT1(16'b0000011100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1900 (
    .a({\picorv32_core/n40 [1],\picorv32_core/n40 [1]}),
    .b({mem_rdata[8],mem_rdata[8]}),
    .c({_al_u1899_o,_al_u1899_o}),
    .d({_al_u1898_o,_al_u1898_o}),
    .mi({open_n10514,_al_u1657_o}),
    .fx({open_n10519,_al_u1900_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~(0*~A))"),
    //.LUTF1("0"),
    //.LUTG0("(~D*~C*~B*~(1*~A))"),
    //.LUTG1("~A*B*~D*C+A*B*~D*C+~A*B*D*C+A*B*D*C"),
    .INIT_LUTF0(16'b0000000000000011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b1100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1901|_al_u2265  (
    .a({open_n10522,_al_u1924_o}),
    .b({_al_u1313_o,_al_u2262_o}),
    .c({\picorv32_core/n667_lutinv ,\picorv32_core/sel41_b0/B5 }),
    .d({open_n10525,\picorv32_core/sel43_b0/B2 }),
    .e({\picorv32_core/pcpi_rs1$0$ ,\picorv32_core/pcpi_rs1$0$ }),
    .f({\picorv32_core/sel43_b0/B2 ,_al_u2265_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(~C*~(0*A)*~(~D*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(~C*~(1*A)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000111100000011),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000010100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1904|picorv32_core/reg15_b32  (
    .a({\picorv32_core/n666_lutinv ,_al_u1902_o}),
    .b({\picorv32_core/n664_lutinv_placeOpt_5 ,\picorv32_core/instr_rdcycleh }),
    .c({\picorv32_core/sel43_b0/B2 ,\picorv32_core/instr_rdinstr }),
    .clk(clk_pad),
    .d({_al_u1903_o,\picorv32_core/count_cycle [32]}),
    .e({\picorv32_core/n543 [0],\picorv32_core/count_instr [0]}),
    .mi({open_n10548,\picorv32_core/n459 [32]}),
    .sr(resetn_placeOpt_8),
    .f({_al_u1904_o,_al_u1903_o}),
    .q({open_n10563,\picorv32_core/count_cycle [32]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~0*~(B*~C)*~(A*~D))"),
    //.LUTF1("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTG0("~(~1*~(B*~C)*~(A*~D))"),
    //.LUTG1("(B*~(~1*~(~A*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110010101110),
    .INIT_LUTF1(16'b0100010000000100),
    .INIT_LUTG0(16'b1111111111111111),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1909|picorv32_core/reg23_b1  (
    .a({\picorv32_core/mem_do_rdata ,_al_u1909_o}),
    .b({\picorv32_core/n669_lutinv_placeOpt_4 ,_al_u1911_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_8 ,_al_u1910_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o,_al_u1908_o}),
    .e({\picorv32_core/mem_wordsize [1],_al_u1912_o}),
    .f({_al_u1909_o,open_n10579}),
    .q({open_n10583,\picorv32_core/mem_wordsize [1]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(~A*~B*~(C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0001000100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1910|picorv32_core/instr_sb_reg  (
    .a({\picorv32_core/mem_do_wdata ,\picorv32_core/is_sb_sh_sw }),
    .b({\picorv32_core/instr_sb ,\picorv32_core/mem_rdata_q [12]}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_8 ,\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({_al_u1546_o,\picorv32_core/mem_rdata_q [14]}),
    .f({_al_u1910_o,open_n10597}),
    .q({open_n10601,\picorv32_core/instr_sb }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~A*B*~(C*~D))"),
    //.LUTF1("(A*~(~0*~(~B*~(C*~D))))"),
    //.LUTG0("(1*~A*B*~(C*~D))"),
    //.LUTG1("(A*~(~1*~(~B*~(C*~D))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0010001000000010),
    .INIT_LUTG0(16'b0100010000000100),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1911|picorv32_core/mem_do_wdata_reg  (
    .a({\picorv32_core/n668_lutinv ,\picorv32_core/mem_do_wdata }),
    .b({\picorv32_core/mem_do_wdata ,\picorv32_core/n668_lutinv }),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_8 ,\picorv32_core/mem_do_prefetch_placeOpt_8 }),
    .ce(\picorv32_core/n747 ),
    .clk(clk_pad),
    .d({_al_u1546_o,_al_u1546_o}),
    .e({\picorv32_core/mem_wordsize [1],resetn_placeOpt_17}),
    .mi({open_n10603,1'b0}),
    .sr(\picorv32_core/n729 ),
    .f({_al_u1911_o,\picorv32_core/n729 }),
    .q({open_n10618,\picorv32_core/mem_do_wdata }));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*A)"),
    //.LUTF1("0"),
    //.LUTG0("(~C*A)"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0000101000001010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000101000001010),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1912|_al_u1609  (
    .a({_al_u1183_o,_al_u1183_o}),
    .c({open_n10621,\picorv32_core/n668_lutinv }),
    .e({\picorv32_core/mem_wordsize [1],open_n10626}),
    .f({_al_u1912_o,_al_u1609_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~0*~(D*~A)*~(C*~B))"),
    //.LUTF1("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTG0("~(~1*~(D*~A)*~(C*~B))"),
    //.LUTG1("(B*~(~1*~(~A*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111010100110000),
    .INIT_LUTF1(16'b0100010000000100),
    .INIT_LUTG0(16'b1111111111111111),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1915|picorv32_core/reg23_b0  (
    .a({\picorv32_core/mem_do_rdata ,_al_u1916_o}),
    .b({\picorv32_core/n669_lutinv_placeOpt_4 ,_al_u1914_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_5 ,_al_u1915_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o_placeOpt_8,_al_u1917_o}),
    .e({\picorv32_core/mem_wordsize [0],_al_u1918_o}),
    .f({_al_u1915_o,open_n10662}),
    .q({open_n10666,\picorv32_core/mem_wordsize [0]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~D*~B*~C*~A+~D*~B*~C*A"),
    //.LUTG0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("~D*~B*~C*~A+~D*~B*C*~A+~D*~B*~C*A+~D*~B*C*A"),
    .INIT_LUTF0(16'b0101010001010100),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0101000001010000),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1916|_al_u1991  (
    .a({open_n10667,\picorv32_core/pcpi_rs1$3$ }),
    .b({\picorv32_core/mem_do_wdata ,\picorv32_core/mem_do_prefetch_placeOpt_5 }),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_5 ,\picorv32_core/mem_do_wdata }),
    .d({\picorv32_core/instr_sh ,open_n10670}),
    .e({_al_u1546_o_placeOpt_8,_al_u1546_o_placeOpt_8}),
    .f({_al_u1916_o,_al_u1991_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUT1("(B*~(~1*~(~A*~(C*~D))))"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b1100110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1917 (
    .a({\picorv32_core/mem_do_wdata ,\picorv32_core/mem_do_wdata }),
    .b({\picorv32_core/n668_lutinv ,\picorv32_core/n668_lutinv }),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_5 ,\picorv32_core/mem_do_prefetch_placeOpt_5 }),
    .d({_al_u1546_o_placeOpt_8,_al_u1546_o_placeOpt_8}),
    .mi({open_n10703,\picorv32_core/mem_wordsize [0]}),
    .fx({open_n10708,_al_u1917_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B*~(C*~D))"),
    //.LUT1("(~B*~A*~(C*~D))"),
    .INIT_LUT0(16'b0001000100000001),
    .INIT_LUT1(16'b0001000100000001),
    .MODE("LOGIC"))
    \_al_u1920|_al_u2225  (
    .a({\picorv32_core/n576 [9],\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_rdata ,\picorv32_core/n576 [12]}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .d({_al_u1546_o_placeOpt_7,_al_u1546_o_placeOpt_7}),
    .f({_al_u1920_o,_al_u2225_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(D*~C)*~(B*~A))"),
    //.LUTF1("(A*~(~0*~(~B*~(C*~D))))"),
    //.LUTG0("~(1*~(D*~C)*~(B*~A))"),
    //.LUTG1("(A*~(~1*~(~B*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0010001000000010),
    .INIT_LUTG0(16'b0100111101000100),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1921|picorv32_core/reg25_b9  (
    .a({\picorv32_core/n669_lutinv_placeOpt_2 ,_al_u1920_o}),
    .b({\picorv32_core/mem_do_rdata ,_al_u1921_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_2 ,_al_u1922_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o_placeOpt_2,_al_u1923_o}),
    .e({\picorv32_core/pcpi_rs1$9$ ,_al_u1932_o}),
    .f({_al_u1921_o,open_n10746}),
    .q({open_n10750,\picorv32_core/pcpi_rs1$9$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(C*~(~1*~B*~(A*~D)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1923 (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .b({\picorv32_core/n576 [9],\picorv32_core/n576 [9]}),
    .c({\picorv32_core/n668_lutinv ,\picorv32_core/n668_lutinv }),
    .d({_al_u1546_o_placeOpt_2,_al_u1546_o_placeOpt_2}),
    .mi({open_n10763,\picorv32_core/mem_do_wdata }),
    .fx({open_n10768,_al_u1923_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1924|_al_u1339  (
    .a({open_n10771,_al_u1338_o}),
    .b({open_n10772,\picorv32_core/n668_lutinv }),
    .c({\picorv32_core/n665_lutinv ,\picorv32_core/n669_lutinv_placeOpt_2 }),
    .d({_al_u1338_o,\picorv32_core/n667_lutinv }),
    .f({_al_u1924_o,_al_u1339_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*~A)"),
    //.LUTF1("(~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*~A)"),
    //.LUTG1("(~B*~A)"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0001000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1926|_al_u1925  (
    .a({_al_u1925_o,\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/decoded_rs1 [1]}),
    .c({open_n10793,\picorv32_core/decoded_rs1 [2]}),
    .d({open_n10796,\picorv32_core/decoded_rs1 [3]}),
    .e({open_n10797,\picorv32_core/decoded_rs1 [4]}),
    .f({_al_u1926_o,_al_u1925_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1100000010100000),
    .MODE("LOGIC"))
    \_al_u1927|_al_u2263  (
    .a({\picorv32_core/cpuregs_p1/dram_do_i0_009 ,_al_u1926_o}),
    .b({\picorv32_core/cpuregs_p1/dram_do_i1_009 ,\picorv32_core/decoded_rs1 [4]}),
    .c({_al_u1926_o,\picorv32_core/cpuregs_p1/dram_do_i0_000 }),
    .d({\picorv32_core/decoded_rs1 [4],\picorv32_core/cpuregs_p1/dram_do_i1_000 }),
    .f({_al_u1927_o,_al_u2263_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(C*~(~A*~(1*B*~D)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010000011100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1928 (
    .a({_al_u1927_o,_al_u1927_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv_placeOpt_4 }),
    .c({\picorv32_core/n664_lutinv_placeOpt_4 ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/instr_lui ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n10850,\picorv32_core/reg_pc [9]}),
    .fx({open_n10855,\picorv32_core/sel41_b9/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*~(B*~D)))"),
    //.LUT1("(~A*~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT_LUT0(16'b0101000001010100),
    .INIT_LUT1(16'b0001000000010101),
    .MODE("LOGIC"))
    \_al_u1929|_al_u1936  (
    .a({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$8$ }),
    .b({\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/mem_do_prefetch_placeOpt_6 }),
    .c({_al_u1302_o,\picorv32_core/mem_do_wdata }),
    .d({\picorv32_core/pcpi_rs1$8$ ,_al_u1546_o_placeOpt_8}),
    .f({_al_u1929_o,_al_u1936_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*A*~B*~C+~D*~A*B*~C+~D*A*B*~C+~D*A*~B*C+~D*~A*B*C+~D*A*B*C"),
    //.LUTF1("A*~D*~C*~B+A*~D*C*~B+A*~D*~C*B+A*~D*C*B"),
    //.LUTG0("~D*~A*B*~C+~D*A*B*~C+~D*~A*B*C+~D*A*B*C"),
    //.LUTG1("A*~D*~C*~B+A*D*~C*~B+A*~D*~C*B+A*D*~C*B"),
    .INIT_LUTF0(16'b0000000011101110),
    .INIT_LUTF1(16'b0000000010101010),
    .INIT_LUTG0(16'b0000000011001100),
    .INIT_LUTG1(16'b0000101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1930|_al_u1969  (
    .a({\picorv32_core/n554 ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .b({open_n10878,\picorv32_core/mem_do_wdata }),
    .c({\picorv32_core/pcpi_rs1$13$ ,open_n10879}),
    .d({\picorv32_core/pcpi_rs1$5$ ,\picorv32_core/pcpi_rs1$5$ }),
    .e({_al_u1302_o,_al_u1546_o_placeOpt_2}),
    .f({_al_u1930_o,_al_u1969_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUTF1("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG0("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0100010001010101),
    .INIT_LUTG0(16'b1010101000000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1932|_al_u1931  (
    .a({\picorv32_core/sel41_b9/B2 ,\picorv32_core/n667_lutinv }),
    .b({_al_u1924_o,_al_u1929_o}),
    .c({open_n10902,_al_u1930_o}),
    .d({\picorv32_core/pcpi_rs1$9$ ,_al_u1313_o}),
    .e({\picorv32_core/sel41_b9/B5 ,\picorv32_core/pcpi_rs1$9$ }),
    .f({_al_u1932_o,\picorv32_core/sel41_b9/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~A*~D*~C*~B+~A*~D*~C*B"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~A*~D*~C*~B+~A*~D*C*~B+~A*~D*~C*B+~A*~D*C*B"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000000000101),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1934|_al_u1937  (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_prefetch_placeOpt_5 }),
    .b({open_n10925,\picorv32_core/n576 [8]}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_5 ,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/n576 [8],_al_u1546_o_placeOpt_8}),
    .e({_al_u1546_o_placeOpt_8,\picorv32_core/mem_do_wdata }),
    .f({_al_u1934_o,_al_u1937_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTF1("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTG0("(B*~(~1*~(~A*~(C*~D))))"),
    //.LUTG1("(B*~(~1*~(~A*~(C*~D))))"),
    .INIT_LUTF0(16'b0100010000000100),
    .INIT_LUTF1(16'b0100010000000100),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1935|_al_u1990  (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/n669_lutinv_placeOpt_3 ,\picorv32_core/n669_lutinv_placeOpt_3 }),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_5 ,\picorv32_core/mem_do_prefetch_placeOpt_5 }),
    .d({_al_u1546_o_placeOpt_5,_al_u1546_o_placeOpt_5}),
    .e({\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/pcpi_rs1$3$ }),
    .f({_al_u1935_o,_al_u1990_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1100000010100000),
    .MODE("LOGIC"))
    \_al_u1938|_al_u2251  (
    .a({\picorv32_core/cpuregs_p1/dram_do_i0_008 ,_al_u1926_o}),
    .b({\picorv32_core/cpuregs_p1/dram_do_i1_008 ,\picorv32_core/decoded_rs1 [4]}),
    .c({_al_u1926_o,\picorv32_core/cpuregs_p1/dram_do_i0_010 }),
    .d({\picorv32_core/decoded_rs1 [4],\picorv32_core/cpuregs_p1/dram_do_i1_010 }),
    .f({_al_u1938_o,_al_u2251_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(D*~(~A*~(1*B*~C)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010111000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1939 (
    .a({_al_u1938_o,_al_u1938_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv_placeOpt_3 }),
    .c({\picorv32_core/instr_lui ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/n664_lutinv_placeOpt_3 ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n11002,\picorv32_core/reg_pc [8]}),
    .fx({open_n11007,\picorv32_core/sel41_b8/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*~(B*~D)))"),
    //.LUT1("(~A*~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT_LUT0(16'b0101000001010100),
    .INIT_LUT1(16'b0000000101010001),
    .MODE("LOGIC"))
    \_al_u1940|_al_u1922  (
    .a({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$9$ }),
    .b({\picorv32_core/pcpi_rs1$7$ ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .c({_al_u1302_o,\picorv32_core/mem_do_wdata }),
    .d({\picorv32_core/pcpi_rs1$9$ ,_al_u1546_o_placeOpt_2}),
    .f({_al_u1940_o,_al_u1922_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*A*~C*~B+~D*~A*C*~B+~D*A*C*~B+~D*A*~C*B+~D*~A*C*B+~D*A*C*B"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+A*B*~C*D+A*B*C*D"),
    //.LUTG0("~D*~A*C*~B+~D*A*C*~B+~D*~A*C*B+~D*A*C*B"),
    //.LUTG1("~A*B*~C*~D+~A*B*C*~D"),
    .INIT_LUTF0(16'b0000000011111010),
    .INIT_LUTF1(16'b1000100011001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1941|_al_u1980  (
    .a({_al_u1302_o,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .b({\picorv32_core/n554 ,open_n11030}),
    .c({open_n11031,\picorv32_core/mem_do_wdata }),
    .d({\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/pcpi_rs1$4$ }),
    .e({\picorv32_core/pcpi_rs1$12$ ,_al_u1546_o_placeOpt_2}),
    .f({_al_u1941_o,_al_u1980_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUTF1("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*A*~D+C*~B*A*~D"),
    //.LUTG0("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    //.LUTG1("~C*~B*A*~D+C*~B*A*~D"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b1010101000000010),
    .INIT_LUTG1(16'b0000000000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1943|_al_u1942  (
    .a({_al_u1924_o,\picorv32_core/n667_lutinv }),
    .b({\picorv32_core/sel41_b8/B5 ,_al_u1940_o}),
    .c({open_n11054,_al_u1941_o}),
    .d({\picorv32_core/sel41_b8/B2 ,_al_u1313_o}),
    .e({\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/pcpi_rs1$8$ }),
    .f({_al_u1943_o,\picorv32_core/sel41_b8/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~C*~B*~D*~A+~C*~B*~D*A"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~C*~B*~D*~A+~C*~B*D*~A+~C*~B*~D*A+~C*~B*D*A"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1945|_al_u1948  (
    .a({open_n11077,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .b({\picorv32_core/n576 [7],\picorv32_core/n576 [7]}),
    .c({\picorv32_core/mem_do_rdata ,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/mem_do_prefetch_placeOpt_2 ,_al_u1546_o_placeOpt_2}),
    .e({_al_u1546_o_placeOpt_2,\picorv32_core/mem_do_wdata }),
    .f({_al_u1945_o,_al_u1948_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(D*~A)*~(B*~C))"),
    //.LUTF1("(A*~(~0*~(~B*~(C*~D))))"),
    //.LUTG0("~(1*~(D*~A)*~(B*~C))"),
    //.LUTG1("(A*~(~1*~(~B*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0010001000000010),
    .INIT_LUTG0(16'b0101110100001100),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1946|picorv32_core/reg25_b7  (
    .a({\picorv32_core/n669_lutinv_placeOpt_2 ,_al_u1947_o}),
    .b({\picorv32_core/mem_do_rdata ,_al_u1946_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_2 ,_al_u1945_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o_placeOpt_2,_al_u1948_o}),
    .e({\picorv32_core/pcpi_rs1$7$ ,_al_u1954_o}),
    .f({_al_u1946_o,open_n11115}),
    .q({open_n11119,\picorv32_core/pcpi_rs1$7$ }));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*D*~C+A*~B*D*C"),
    //.LUTF1("A*~B*D*~C+A*~B*D*C"),
    //.LUTG0("A*B*~D*~C+A*~B*D*~C+A*B*D*~C+A*B*~D*C+A*~B*D*C+A*B*D*C"),
    //.LUTG1("A*B*~D*~C+A*~B*D*~C+A*B*D*~C+A*B*~D*C+A*~B*D*C+A*B*D*C"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0010001000000000),
    .INIT_LUTG0(16'b1010101010001000),
    .INIT_LUTG1(16'b1010101010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1949|_al_u2240  (
    .a({_al_u1926_o,_al_u1926_o}),
    .b({\picorv32_core/decoded_rs1 [4],\picorv32_core/decoded_rs1 [4]}),
    .d({\picorv32_core/cpuregs_p1/dram_do_i0_007 ,\picorv32_core/cpuregs_p1/dram_do_i0_011 }),
    .e({\picorv32_core/cpuregs_p1/dram_do_i1_007 ,\picorv32_core/cpuregs_p1/dram_do_i1_011 }),
    .f({_al_u1949_o,_al_u2240_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*~(B*~D)))"),
    //.LUT1("(~A*~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT_LUT0(16'b0101000001010100),
    .INIT_LUT1(16'b0000000101010001),
    .MODE("LOGIC"))
    \_al_u1951|_al_u1958  (
    .a({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$6$ }),
    .b({\picorv32_core/pcpi_rs1$6$ ,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .c({_al_u1302_o,\picorv32_core/mem_do_wdata }),
    .d({\picorv32_core/pcpi_rs1$8$ ,_al_u1546_o_placeOpt_7}),
    .f({_al_u1951_o,_al_u1958_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUT1("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1953 (
    .a({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .b({_al_u1951_o,_al_u1951_o}),
    .c({_al_u1952_o,_al_u1952_o}),
    .d({_al_u1313_o,_al_u1313_o}),
    .mi({open_n11176,\picorv32_core/pcpi_rs1$7$ }),
    .fx({open_n11181,\picorv32_core/sel41_b7/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("~A*~B*~D*~C+~A*~B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("~A*~B*D*~C+~A*~B*D*C"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0001000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1954|_al_u1950  (
    .a({\picorv32_core/sel41_b7/B5 ,_al_u1949_o}),
    .b({\picorv32_core/sel41_b7/B2 ,\picorv32_core/n664_lutinv_placeOpt_2 }),
    .c({open_n11184,\picorv32_core/instr_lui }),
    .d({_al_u1924_o,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/pcpi_rs1$7$ ,\picorv32_core/reg_pc [7]}),
    .f({_al_u1954_o,\picorv32_core/sel41_b7/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B*~(C*~D))"),
    //.LUT1("(~B*~A*~(C*~D))"),
    .INIT_LUT0(16'b0001000100000001),
    .INIT_LUT1(16'b0001000100000001),
    .MODE("LOGIC"))
    \_al_u1956|_al_u2214  (
    .a({\picorv32_core/n576 [6],\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_rdata ,\picorv32_core/n576 [13]}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_7 ,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .d({_al_u1546_o_placeOpt_7,_al_u1546_o_placeOpt_7}),
    .f({_al_u1956_o,_al_u2214_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(A*~C)*~(D*~B))"),
    //.LUTF1("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTG0("~(1*~(A*~C)*~(D*~B))"),
    //.LUTG1("(B*~(~1*~(~A*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0100010000000100),
    .INIT_LUTG0(16'b0011101100001010),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1957|picorv32_core/reg25_b6  (
    .a({\picorv32_core/mem_do_rdata ,_al_u1959_o}),
    .b({\picorv32_core/n669_lutinv_placeOpt_2 ,_al_u1956_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_7 ,_al_u1958_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o_placeOpt_7,_al_u1957_o}),
    .e({\picorv32_core/pcpi_rs1$6$ ,_al_u1965_o}),
    .f({_al_u1957_o,open_n11242}),
    .q({open_n11246,\picorv32_core/pcpi_rs1$6$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(A*~(~1*~B*~(D*~C)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1959 (
    .a({\picorv32_core/n668_lutinv ,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .b({\picorv32_core/n576 [6],\picorv32_core/n576 [6]}),
    .c({_al_u1546_o_placeOpt_1,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/mem_do_prefetch_placeOpt_7 ,_al_u1546_o_placeOpt_1}),
    .mi({open_n11259,\picorv32_core/mem_do_wdata }),
    .fx({open_n11264,_al_u1959_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*C*~D+A*~B*C*D"),
    //.LUTF1("A*~B*D*~C+A*~B*D*C"),
    //.LUTG0("A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG1("A*B*~D*~C+A*~B*D*~C+A*B*D*~C+A*B*~D*C+A*~B*D*C+A*B*D*C"),
    .INIT_LUTF0(16'b0010000000100000),
    .INIT_LUTF1(16'b0010001000000000),
    .INIT_LUTG0(16'b1010100010101000),
    .INIT_LUTG1(16'b1010101010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1960|_al_u2229  (
    .a({_al_u1926_o,_al_u1926_o}),
    .b({\picorv32_core/decoded_rs1 [4],\picorv32_core/decoded_rs1 [4]}),
    .c({open_n11267,\picorv32_core/cpuregs_p1/dram_do_i0_012 }),
    .d({\picorv32_core/cpuregs_p1/dram_do_i0_006 ,open_n11270}),
    .e({\picorv32_core/cpuregs_p1/dram_do_i1_006 ,\picorv32_core/cpuregs_p1/dram_do_i1_012 }),
    .f({_al_u1960_o,_al_u2229_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*((~C*~A)*~(0)*~(D)+(~C*~A)*0*~(D)+~((~C*~A))*0*D+(~C*~A)*0*D))"),
    //.LUTF1("~A*~D*~C*~B+~A*~D*C*~B+~A*D*C*~B+~A*~D*~C*B+~A*~D*C*B+~A*D*C*B"),
    //.LUTG0("(B*((~C*~A)*~(1)*~(D)+(~C*~A)*1*~(D)+~((~C*~A))*1*D+(~C*~A)*1*D))"),
    //.LUTG1("~A*~D*~C*~B+~A*~D*~C*B"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b0101000001010101),
    .INIT_LUTG0(16'b1100110000000100),
    .INIT_LUTG1(16'b0000000000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1962|_al_u1964  (
    .a({\picorv32_core/n554 ,_al_u1962_o}),
    .b({open_n11291,\picorv32_core/n667_lutinv }),
    .c({_al_u1302_o,_al_u1963_o}),
    .d({\picorv32_core/pcpi_rs1$5$ ,_al_u1313_o}),
    .e({\picorv32_core/pcpi_rs1$7$ ,\picorv32_core/pcpi_rs1$6$ }),
    .f({_al_u1962_o,\picorv32_core/sel41_b6/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0000000011011101),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1965|_al_u1961  (
    .a({\picorv32_core/pcpi_rs1$6$ ,_al_u1960_o}),
    .b({_al_u1924_o,\picorv32_core/n664_lutinv_placeOpt_2 }),
    .c({open_n11314,\picorv32_core/instr_lui }),
    .d({\picorv32_core/sel41_b6/B5 ,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/sel41_b6/B2 ,\picorv32_core/reg_pc [6]}),
    .f({_al_u1965_o,\picorv32_core/sel41_b6/B5 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+~A*C*B*D"),
    //.LUTF1("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("0"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0101010100010001),
    .INIT_LUTF1(16'b0101010100010001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1967|_al_u2181  (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .d({_al_u1546_o_placeOpt_2,_al_u1546_o_placeOpt_2}),
    .e({\picorv32_core/n576 [5],\picorv32_core/n576 [16]}),
    .f({_al_u1967_o,_al_u2181_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUT1("(C*~(~1*~(~A*~(B*~D))))"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b1111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1968 (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/n669_lutinv_placeOpt_2 }),
    .c({\picorv32_core/n669_lutinv_placeOpt_2 ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .d({_al_u1546_o_placeOpt_2,_al_u1546_o_placeOpt_2}),
    .mi({open_n11373,\picorv32_core/pcpi_rs1$5$ }),
    .fx({open_n11378,_al_u1968_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(C*~(~1*~B*~(A*~D)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1970 (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .b({\picorv32_core/n576 [5],\picorv32_core/n576 [5]}),
    .c({\picorv32_core/n668_lutinv ,\picorv32_core/n668_lutinv }),
    .d({_al_u1546_o_placeOpt_2,_al_u1546_o_placeOpt_2}),
    .mi({open_n11393,\picorv32_core/mem_do_wdata }),
    .fx({open_n11398,_al_u1970_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010110000000000),
    .MODE("LOGIC"))
    \_al_u1971|_al_u2218  (
    .a({\picorv32_core/cpuregs_p1/dram_do_i1_005 ,_al_u1926_o}),
    .b({\picorv32_core/cpuregs_p1/dram_do_i0_005 ,\picorv32_core/decoded_rs1 [4]}),
    .c({\picorv32_core/decoded_rs1 [4],\picorv32_core/cpuregs_p1/dram_do_i0_013 }),
    .d({_al_u1926_o,\picorv32_core/cpuregs_p1/dram_do_i1_013 }),
    .f({_al_u1971_o,_al_u2218_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(C*~(~A*~(1*B*~D)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010000011100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1972 (
    .a({_al_u1971_o,_al_u1971_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv }),
    .c({\picorv32_core/n664_lutinv ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/instr_lui ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n11433,\picorv32_core/reg_pc [5]}),
    .fx({open_n11438,\picorv32_core/sel41_b5/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUT1("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1975 (
    .a({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .b({_al_u1973_o,_al_u1973_o}),
    .c({_al_u1974_o,_al_u1974_o}),
    .d({_al_u1313_o,_al_u1313_o}),
    .mi({open_n11453,\picorv32_core/pcpi_rs1$5$ }),
    .fx({open_n11458,\picorv32_core/sel41_b5/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+~A*B*~C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*B*C*D"),
    //.LUTF1("~C*~B*~A*~D+~C*~B*A*~D+~C*~B*~A*D+~C*B*~A*D+~C*~B*A*D+~C*B*A*D"),
    //.LUTG0("~A*~B*~C*~D+~A*~B*~C*D"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0100010101000101),
    .INIT_LUTF1(16'b0000111100000011),
    .INIT_LUTG0(16'b0000000100000001),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1976|_al_u1984  (
    .a({open_n11461,\picorv32_core/n554 }),
    .b({\picorv32_core/pcpi_rs1$5$ ,_al_u1302_o}),
    .c({\picorv32_core/sel41_b5/B5 ,\picorv32_core/pcpi_rs1$3$ }),
    .d({_al_u1924_o,open_n11464}),
    .e({\picorv32_core/sel41_b5/B2 ,\picorv32_core/pcpi_rs1$5$ }),
    .f({_al_u1976_o,_al_u1984_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~A*~D*~B*~C+~A*~D*~B*C"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~A*~D*~B*~C+~A*~D*B*~C+~A*~D*~B*C+~A*~D*B*C"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000000010001),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1978|_al_u1981  (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/n576 [4]}),
    .c({open_n11485,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/n576 [4],_al_u1546_o_placeOpt_2}),
    .e({_al_u1546_o_placeOpt_2,\picorv32_core/mem_do_wdata }),
    .f({_al_u1978_o,_al_u1981_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(C*~B)*~(D*~A))"),
    //.LUTF1("(A*~(~0*~(~B*~(C*~D))))"),
    //.LUTG0("~(1*~(C*~B)*~(D*~A))"),
    //.LUTG1("(A*~(~1*~(~B*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0010001000000010),
    .INIT_LUTG0(16'b0111010100110000),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1979|picorv32_core/reg25_b4  (
    .a({\picorv32_core/n669_lutinv_placeOpt_2 ,_al_u1978_o}),
    .b({\picorv32_core/mem_do_rdata ,_al_u1980_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_2 ,_al_u1981_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o_placeOpt_2,_al_u1979_o}),
    .e({\picorv32_core/pcpi_rs1$4$ ,_al_u1987_o}),
    .f({_al_u1979_o,open_n11523}),
    .q({open_n11527,\picorv32_core/pcpi_rs1$4$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1100000010100000),
    .MODE("LOGIC"))
    \_al_u1982|_al_u2207  (
    .a({\picorv32_core/cpuregs_p1/dram_do_i0_004 ,_al_u1926_o}),
    .b({\picorv32_core/cpuregs_p1/dram_do_i1_004 ,\picorv32_core/decoded_rs1 [4]}),
    .c({_al_u1926_o,\picorv32_core/cpuregs_p1/dram_do_i0_014 }),
    .d({\picorv32_core/decoded_rs1 [4],\picorv32_core/cpuregs_p1/dram_do_i1_014 }),
    .f({_al_u1982_o,_al_u2207_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~D*~(0*A*~C)))"),
    //.LUT1("(A*~(~D*~(1*B*~C)))"),
    .INIT_LUT0(16'b1100110000000000),
    .INIT_LUT1(16'b1010101000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1983 (
    .a({\picorv32_core/n664_lutinv ,\picorv32_core/is_lui_auipc_jal }),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv }),
    .c({\picorv32_core/instr_lui ,\picorv32_core/instr_lui }),
    .d({_al_u1982_o,_al_u1982_o}),
    .mi({open_n11560,\picorv32_core/reg_pc [4]}),
    .fx({open_n11565,\picorv32_core/sel41_b4/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUT1("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1986 (
    .a({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .b({_al_u1984_o,_al_u1984_o}),
    .c({_al_u1985_o,_al_u1985_o}),
    .d({_al_u1313_o,_al_u1313_o}),
    .mi({open_n11580,\picorv32_core/pcpi_rs1$4$ }),
    .fx({open_n11585,\picorv32_core/sel41_b4/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*~C*~A+~B*D*~C*~A+~B*D*C*~A+~B*~D*~C*A+~B*D*~C*A+~B*D*C*A"),
    //.LUTF1("~A*~B*~D*~C+~A*~B*D*~C+~A*B*D*~C+~A*~B*~D*C+~A*~B*D*C+~A*B*D*C"),
    //.LUTG0("~B*~D*~C*~A+~B*~D*~C*A"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b0101010100010001),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1987|_al_u1973  (
    .a({\picorv32_core/sel41_b4/B2 ,open_n11588}),
    .b({\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/n554 }),
    .c({open_n11589,\picorv32_core/pcpi_rs1$4$ }),
    .d({_al_u1924_o,_al_u1302_o}),
    .e({\picorv32_core/sel41_b4/B5 ,\picorv32_core/pcpi_rs1$6$ }),
    .f({_al_u1987_o,_al_u1973_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~A*~D*~B*~C+~A*~D*~B*C"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~A*~D*~B*~C+~A*~D*B*~C+~A*~D*~B*C+~A*~D*B*C"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000000010001),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1989|_al_u1992  (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_prefetch_placeOpt_5 }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_5 ,\picorv32_core/n576 [3]}),
    .c({open_n11612,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/n576 [3],_al_u1546_o_placeOpt_5}),
    .e({_al_u1546_o_placeOpt_5,\picorv32_core/mem_do_wdata }),
    .f({_al_u1989_o,_al_u1992_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*C*~D+A*B*C*~D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("A*~D*C*~B+A*~D*C*B"),
    //.LUTG0("A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG1("A*D*~C*~B+A*~D*C*~B+A*D*C*~B+A*D*~C*B+A*~D*C*B+A*D*C*B"),
    .INIT_LUTF0(16'b1010000010100000),
    .INIT_LUTF1(16'b0000000010100000),
    .INIT_LUTG0(16'b1010101000000000),
    .INIT_LUTG1(16'b1010101010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1993|_al_u2196  (
    .a({_al_u1926_o,_al_u1926_o}),
    .c({\picorv32_core/cpuregs_p1/dram_do_i0_003 ,\picorv32_core/cpuregs_p1/dram_do_i0_015 }),
    .d({\picorv32_core/decoded_rs1 [4],\picorv32_core/cpuregs_p1/dram_do_i1_015 }),
    .e({\picorv32_core/cpuregs_p1/dram_do_i1_003 ,\picorv32_core/decoded_rs1 [4]}),
    .f({_al_u1993_o,_al_u2196_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+~(A)*B*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+A*B*~(C)*D*~(0)+A*~(B)*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(D)*~(C)*~(B)*~(1)+A*~(D)*~(C)*~(B)*~(1)+~(A)*D*~(C)*~(B)*~(1)+A*D*~(C)*~(B)*~(1)+A*~(D)*C*~(B)*~(1)+~(A)*D*C*~(B)*~(1)+A*D*C*~(B)*~(1)+~(A)*~(D)*~(C)*B*~(1)+A*~(D)*~(C)*B*~(1)+A*D*~(C)*B*~(1)+A*~(D)*C*B*~(1)+A*D*C*B*~(1)+~(A)*~(D)*~(C)*~(B)*1+A*~(D)*~(C)*~(B)*1+~(A)*D*~(C)*~(B)*1+A*~(D)*C*~(B)*1+~(A)*D*C*~(B)*1+~(A)*~(D)*~(C)*B*1+A*~(D)*~(C)*B*1+A*~(D)*C*B*1)"),
    .INIT_LUT0(16'b1010101111101111),
    .INIT_LUT1(16'b0001000110101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1995 (
    .a({\picorv32_core/n554 ,\picorv32_core/n554 }),
    .b({\picorv32_core/pcpi_rs1$4$ ,_al_u1302_o}),
    .c({\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$2$ }),
    .d({_al_u1302_o,\picorv32_core/pcpi_rs1$4$ }),
    .mi({open_n11671,\picorv32_core/pcpi_rs1$7$ }),
    .fx({open_n11676,_al_u1995_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("(~D*~(B*(~C*~(0)*~(A)+~C*0*~(A)+~(~C)*0*A+~C*0*A)))"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("(~D*~(B*(~C*~(1)*~(A)+~C*1*~(A)+~(~C)*1*A+~C*1*A)))"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0000000011111011),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0000000001110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1996|_al_u1994  (
    .a({_al_u1313_o,_al_u1993_o}),
    .b({\picorv32_core/n667_lutinv ,\picorv32_core/n664_lutinv_placeOpt_2 }),
    .c({_al_u1995_o,\picorv32_core/instr_lui }),
    .d({\picorv32_core/sel41_b3/B5 ,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/pcpi_rs1$3$ ,\picorv32_core/reg_pc [3]}),
    .f({_al_u1996_o,\picorv32_core/sel41_b3/B5 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    //.LUTF1("~A*~B*~D*~C+~A*~B*~D*C"),
    //.LUTG0("~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG1("~A*~B*~D*~C+~A*B*~D*~C+~A*~B*~D*C+~A*B*~D*C"),
    .INIT_LUTF0(16'b0001000100010001),
    .INIT_LUTF1(16'b0000000000010001),
    .INIT_LUTG0(16'b0001000100000000),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1999|_al_u2170  (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_6 ,\picorv32_core/n576 [17]}),
    .d({\picorv32_core/n576 [31],_al_u1546_o_placeOpt_6}),
    .e({_al_u1546_o_placeOpt_6,\picorv32_core/mem_do_prefetch_placeOpt_6 }),
    .f({_al_u1999_o,_al_u2170_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTF1("A*~D*~C*~B+~A*~D*C*~B+A*~D*C*~B+A*~D*~C*B+~A*~D*C*B+A*~D*C*B"),
    //.LUTG0("(B*~(~1*~(~A*~(C*~D))))"),
    //.LUTG1("~A*~D*C*~B+A*~D*C*~B+~A*~D*C*B+A*~D*C*B"),
    .INIT_LUTF0(16'b0100010000000100),
    .INIT_LUTF1(16'b0000000011111010),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2001|_al_u2000  (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_6 ,\picorv32_core/mem_do_rdata }),
    .b({open_n11725,\picorv32_core/n669_lutinv_placeOpt_3 }),
    .c({\picorv32_core/mem_do_wdata ,\picorv32_core/mem_do_prefetch_placeOpt_6 }),
    .d({\picorv32_core/pcpi_rs1$31$ ,_al_u1546_o_placeOpt_6}),
    .e({_al_u1546_o_placeOpt_6,\picorv32_core/pcpi_rs1$31$ }),
    .f({_al_u2001_o,_al_u2000_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(A*~(~1*~B*~(C*~D)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2002 (
    .a({\picorv32_core/n668_lutinv ,\picorv32_core/mem_do_prefetch_placeOpt_6 }),
    .b({\picorv32_core/n576 [31],\picorv32_core/n576 [31]}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_6 ,\picorv32_core/n668_lutinv }),
    .d({_al_u1546_o_placeOpt_6,_al_u1546_o_placeOpt_6}),
    .mi({open_n11760,\picorv32_core/mem_do_wdata }),
    .fx({open_n11765,_al_u2002_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("0"),
    //.LUTG0("~C*~B*A*~D+C*~B*A*~D+~C*B*~A*D+C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG1("~C*~B*D*~A+C*~B*D*~A+~C*B*~D*A+C*B*~D*A+~C*~B*D*A+C*~B*D*A+~C*B*D*A+C*B*D*A"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1110111000100010),
    .INIT_LUTG1(16'b1011101110001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2003|_al_u2185  (
    .a({\picorv32_core/cpuregs_p1/dram_do_i1_031 ,\picorv32_core/cpuregs_p1/dram_do_i0_016 }),
    .b({\picorv32_core/decoded_rs1 [4],\picorv32_core/decoded_rs1 [4]}),
    .d({\picorv32_core/cpuregs_p1/dram_do_i0_031 ,\picorv32_core/cpuregs_p1/dram_do_i1_016 }),
    .e({_al_u1926_o,_al_u1926_o}),
    .f({_al_u2003_o,_al_u2185_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b0000000011100100),
    .MODE("LOGIC"))
    \_al_u2005|_al_u2044  (
    .a({\picorv32_core/n554 ,\picorv32_core/n554 }),
    .b({\picorv32_core/pcpi_rs1$30$ ,_al_u1302_o}),
    .c({\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/pcpi_rs1$27$ }),
    .d({_al_u1302_o,\picorv32_core/pcpi_rs1$29$ }),
    .f({_al_u2005_o,_al_u2044_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("(~A*~(D*B)*~(0*~C))"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("(~A*~(D*B)*~(1*~C))"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0001000101010101),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2007|_al_u2004  (
    .a({\picorv32_core/sel41_b31/B5 ,_al_u2003_o}),
    .b({\picorv32_core/n570 [31],\picorv32_core/n664_lutinv_placeOpt_2 }),
    .c({_al_u1924_o,\picorv32_core/instr_lui }),
    .d({\picorv32_core/n667_lutinv ,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/pcpi_rs1$31$ ,\picorv32_core/reg_pc [31]}),
    .f({_al_u2007_o,\picorv32_core/sel41_b31/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B*~(C*~D))"),
    //.LUT1("(~B*~A*~(C*~D))"),
    .INIT_LUT0(16'b0001000100000001),
    .INIT_LUT1(16'b0001000100000001),
    .MODE("LOGIC"))
    \_al_u2009|_al_u2138  (
    .a({\picorv32_core/n576 [30],\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_rdata ,\picorv32_core/n576 [1]}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_7 ,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .d({_al_u1546_o_placeOpt_7,_al_u1546_o_placeOpt_7}),
    .f({_al_u2009_o,_al_u2138_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(D*~A)*~(B*~C))"),
    //.LUTF1("(A*~(~0*~(~B*~(C*~D))))"),
    //.LUTG0("~(1*~(D*~A)*~(B*~C))"),
    //.LUTG1("(A*~(~1*~(~B*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0010001000000010),
    .INIT_LUTG0(16'b0101110100001100),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2010|picorv32_core/reg25_b30  (
    .a({\picorv32_core/n669_lutinv_placeOpt_2 ,_al_u2011_o}),
    .b({\picorv32_core/mem_do_rdata ,_al_u2010_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_7 ,_al_u2009_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o_placeOpt_7,_al_u2012_o}),
    .e({\picorv32_core/pcpi_rs1$30$ ,_al_u2018_o}),
    .f({_al_u2010_o,open_n11869}),
    .q({open_n11873,\picorv32_core/pcpi_rs1$30$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(A*~(~1*~B*~(D*~C)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2012 (
    .a({\picorv32_core/n668_lutinv ,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .b({\picorv32_core/n576 [30],\picorv32_core/n576 [30]}),
    .c({_al_u1546_o_placeOpt_7,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/mem_do_prefetch_placeOpt_7 ,_al_u1546_o_placeOpt_7}),
    .mi({open_n11886,\picorv32_core/mem_do_wdata }),
    .fx({open_n11891,_al_u2012_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*B*~(C*~(0*~D)))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*B*C*D"),
    //.LUTG0("(~A*B*~(C*~(1*~D)))"),
    //.LUTG1("~A*~B*~C*~D+~A*~B*~C*D"),
    .INIT_LUTF0(16'b0000010000000100),
    .INIT_LUTF1(16'b0100010101000101),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2013|_al_u2015  (
    .a({\picorv32_core/n554 ,_al_u2013_o}),
    .b({_al_u1302_o,\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv }),
    .c({\picorv32_core/pcpi_rs1$29$ ,_al_u2014_o}),
    .d({open_n11896,_al_u1302_o}),
    .e({\picorv32_core/pcpi_rs1$31$ ,\picorv32_core/pcpi_rs1$26$ }),
    .f({_al_u2013_o,_al_u2015_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B)*~((~D*~C))*~(0)+A*~(B)*(~D*~C)*~(0)+~(A)*~(B)*~((~D*~C))*0+A*~(B)*~((~D*~C))*0+~(A)*B*~((~D*~C))*0+A*B*~((~D*~C))*0+A*~(B)*(~D*~C)*0+~(A)*B*(~D*~C)*0+A*B*(~D*~C)*0)"),
    //.LUTF1("C*~B*~A*~D+C*B*~A*~D+C*~B*A*~D+C*B*A*~D+C*~B*~A*D+C*~B*A*D"),
    //.LUTG0("(A*~(B)*~((~D*~C))*~(1)+A*~(B)*(~D*~C)*~(1)+~(A)*~(B)*~((~D*~C))*1+A*~(B)*~((~D*~C))*1+~(A)*B*~((~D*~C))*1+A*B*~((~D*~C))*1+A*~(B)*(~D*~C)*1+~(A)*B*(~D*~C)*1+A*B*(~D*~C)*1)"),
    //.LUTG1("C*~B*~A*~D+C*B*~A*~D+C*~B*A*~D+C*B*A*~D"),
    .INIT_LUTF0(16'b0010001000100010),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b1111111111111110),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2014|_al_u2006  (
    .a({open_n11917,_al_u2005_o}),
    .b({\picorv32_core/instr_sra ,_al_u1313_o}),
    .c({\picorv32_core/n554 ,\picorv32_core/instr_sra }),
    .d({\picorv32_core/pcpi_rs1$31$ ,\picorv32_core/instr_srai }),
    .e({\picorv32_core/instr_srai ,\picorv32_core/pcpi_rs1$31$ }),
    .f({_al_u2014_o,\picorv32_core/n570 [31]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010110000000000),
    .MODE("LOGIC"))
    \_al_u2016|_al_u2174  (
    .a({\picorv32_core/cpuregs_p1/dram_do_i1_030 ,_al_u1926_o}),
    .b({\picorv32_core/cpuregs_p1/dram_do_i0_030 ,\picorv32_core/decoded_rs1 [4]}),
    .c({\picorv32_core/decoded_rs1 [4],\picorv32_core/cpuregs_p1/dram_do_i0_017 }),
    .d({_al_u1926_o,\picorv32_core/cpuregs_p1/dram_do_i1_017 }),
    .f({_al_u2016_o,_al_u2174_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(C*~(~A*~(1*B*~D)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010000011100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2017 (
    .a({_al_u2016_o,_al_u2016_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv }),
    .c({\picorv32_core/n664_lutinv ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/instr_lui ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n11972,\picorv32_core/reg_pc [30]}),
    .fx({open_n11977,\picorv32_core/sel41_b30/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*~(0*~A))"),
    //.LUT1("(~D*~C*~B*~(1*~A))"),
    .INIT_LUT0(16'b0000000000000011),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2018 (
    .a({_al_u1924_o,_al_u1924_o}),
    .b({_al_u2015_o,_al_u2015_o}),
    .c({\picorv32_core/sel41_b30/B5 ,\picorv32_core/sel41_b30/B5 }),
    .d({\picorv32_core/sel43_b30/B2 ,\picorv32_core/sel43_b30/B2 }),
    .mi({open_n11992,\picorv32_core/pcpi_rs1$30$ }),
    .fx({open_n11997,_al_u2018_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~A*~B*~C*~D+~A*~B*~C*D"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000100000001),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0001000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2020|_al_u2023  (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .b({\picorv32_core/n576 [2],\picorv32_core/n576 [2]}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/n668_lutinv }),
    .d({open_n12002,_al_u1546_o_placeOpt_2}),
    .e({_al_u1546_o_placeOpt_2,\picorv32_core/mem_do_wdata }),
    .f({_al_u2020_o,_al_u2023_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTF1("~D*B*~A*~C+~D*~B*A*~C+~D*B*A*~C+~D*B*~A*C+~D*~B*A*C+~D*B*A*C"),
    //.LUTG0("(B*~(~1*~(~A*~(C*~D))))"),
    //.LUTG1("~D*~B*A*~C+~D*B*A*~C+~D*~B*A*C+~D*B*A*C"),
    .INIT_LUTF0(16'b0100010000000100),
    .INIT_LUTF1(16'b0000000011101110),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b0000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2022|_al_u2021  (
    .a({\picorv32_core/mem_do_wdata ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/n669_lutinv_placeOpt_2 }),
    .c({open_n12023,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .d({\picorv32_core/pcpi_rs1$2$ ,_al_u1546_o_placeOpt_2}),
    .e({_al_u1546_o_placeOpt_2,\picorv32_core/pcpi_rs1$2$ }),
    .f({_al_u2022_o,_al_u2021_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010110000000000),
    .MODE("LOGIC"))
    \_al_u2024|_al_u2163  (
    .a({\picorv32_core/cpuregs_p1/dram_do_i1_002 ,_al_u1926_o}),
    .b({\picorv32_core/cpuregs_p1/dram_do_i0_002 ,\picorv32_core/decoded_rs1 [4]}),
    .c({\picorv32_core/decoded_rs1 [4],\picorv32_core/cpuregs_p1/dram_do_i0_018 }),
    .d({_al_u1926_o,\picorv32_core/cpuregs_p1/dram_do_i1_018 }),
    .f({_al_u2024_o,_al_u2163_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(C*~(~A*~(1*B*~D)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010000011100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2025 (
    .a({_al_u2024_o,_al_u2024_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv }),
    .c({\picorv32_core/n664_lutinv ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/instr_lui ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n12078,\picorv32_core/reg_pc [2]}),
    .fx({open_n12083,\picorv32_core/sel41_b2/B5 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+~(A)*B*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+A*B*~(C)*D*~(0)+A*~(B)*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("(~A*~(B*(~D*~(0)*~(C)+~D*0*~(C)+~(~D)*0*C+~D*0*C)))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+~(A)*B*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+A*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+A*B*~(C)*D*~(1)+A*~(B)*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("(~A*~(B*(~D*~(1)*~(C)+~D*1*~(C)+~(~D)*1*C+~D*1*C)))"),
    .INIT_LUTF0(16'b1010101111101111),
    .INIT_LUTF1(16'b0101010101010001),
    .INIT_LUTG0(16'b0010001101100111),
    .INIT_LUTG1(16'b0001010100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2027|_al_u2026  (
    .a({\picorv32_core/sel41_b2/B5 ,\picorv32_core/n554 }),
    .b({\picorv32_core/n667_lutinv ,_al_u1302_o}),
    .c({_al_u1313_o,\picorv32_core/pcpi_rs1$1$ }),
    .d({_al_u2026_o,\picorv32_core/pcpi_rs1$3$ }),
    .e({\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$6$ }),
    .f({_al_u2027_o,_al_u2026_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*B*D)"),
    //.LUT1("(D*~(B*~A))"),
    .INIT_LUT0(16'b1000100000000000),
    .INIT_LUT1(16'b1011101100000000),
    .MODE("LOGIC"))
    \_al_u2028|_al_u1724  (
    .a({_al_u1924_o,\picorv32_core/pcpi_rs1$30$ }),
    .b({\picorv32_core/pcpi_rs1$2$ ,_al_u1313_o}),
    .d({_al_u2027_o,\picorv32_core/n667_lutinv }),
    .f({_al_u2028_o,\picorv32_core/sel43_b30/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~D*~B*~C*~A+~D*~B*~C*A"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~D*~B*~C*~A+~D*~B*C*~A+~D*~B*~C*A+~D*~B*C*A"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2030|_al_u2033  (
    .a({open_n12130,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .b({\picorv32_core/n576 [29],\picorv32_core/n576 [29]}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_7 ,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/mem_do_rdata ,_al_u1546_o_placeOpt_7}),
    .e({_al_u1546_o_placeOpt_7,\picorv32_core/mem_do_wdata }),
    .f({_al_u2030_o,_al_u2033_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(C*~B)*~(A*~D))"),
    //.LUTF1("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTG0("~(1*~(C*~B)*~(A*~D))"),
    //.LUTG1("(B*~(~1*~(~A*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0100010000000100),
    .INIT_LUTG0(16'b0011000010111010),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2031|picorv32_core/reg25_b29  (
    .a({\picorv32_core/mem_do_rdata ,_al_u2031_o}),
    .b({\picorv32_core/n669_lutinv_placeOpt_2 ,_al_u2032_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_2 ,_al_u2033_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o_placeOpt_2,_al_u2030_o}),
    .e({\picorv32_core/pcpi_rs1$29$ ,_al_u2038_o}),
    .f({_al_u2031_o,open_n12168}),
    .q({open_n12172,\picorv32_core/pcpi_rs1$29$ }));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*C*~(B*~(0*~D)))"),
    //.LUTF1("~C*~B*~A*~D+~C*B*~A*~D+~C*~B*A*~D+~C*B*A*~D+~C*~B*~A*D+~C*~B*A*D"),
    //.LUTG0("(~A*C*~(B*~(1*~D)))"),
    //.LUTG1("~C*B*~A*~D+~C*B*A*~D"),
    .INIT_LUTF0(16'b0001000000010000),
    .INIT_LUTF1(16'b0000001100001111),
    .INIT_LUTG0(16'b0001000001010000),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2034|_al_u2035  (
    .a({open_n12173,_al_u2034_o}),
    .b({_al_u1302_o,_al_u2014_o}),
    .c({\picorv32_core/n554 ,\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv }),
    .d({\picorv32_core/pcpi_rs1$30$ ,_al_u1302_o}),
    .e({\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/pcpi_rs1$25$ }),
    .f({_al_u2034_o,_al_u2035_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("0"),
    //.LUTG0("~C*~B*D*~A+C*~B*D*~A+~C*B*~D*A+C*B*~D*A+~C*~B*D*A+C*~B*D*A+~C*B*D*A+C*B*D*A"),
    //.LUTG1("~D*~B*C*~A+D*~B*C*~A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1011101110001000),
    .INIT_LUTG1(16'b1011100010111000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2036|_al_u2152  (
    .a({\picorv32_core/cpuregs_p1/dram_do_i1_029 ,\picorv32_core/cpuregs_p1/dram_do_i1_019 }),
    .b({\picorv32_core/decoded_rs1 [4],\picorv32_core/decoded_rs1 [4]}),
    .c({\picorv32_core/cpuregs_p1/dram_do_i0_029 ,open_n12196}),
    .d({open_n12199,\picorv32_core/cpuregs_p1/dram_do_i0_019 }),
    .e({_al_u1926_o,_al_u1926_o}),
    .f({_al_u2036_o,_al_u2152_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("(~D*~A*~B*~(0*~C))"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("(~D*~A*~B*~(1*~C))"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0000000000010001),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0000000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2038|_al_u2037  (
    .a({\picorv32_core/sel41_b29/B5 ,_al_u2036_o}),
    .b({_al_u2035_o,\picorv32_core/n664_lutinv_placeOpt_1 }),
    .c({_al_u1924_o,\picorv32_core/instr_lui }),
    .d({\picorv32_core/sel43_b29/B2 ,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/pcpi_rs1$29$ ,\picorv32_core/reg_pc [29]}),
    .f({_al_u2038_o,\picorv32_core/sel41_b29/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B*~(C*~D))"),
    //.LUT1("(~C*~B*~(A*~D))"),
    .INIT_LUT0(16'b0001000100000001),
    .INIT_LUT1(16'b0000001100000001),
    .MODE("LOGIC"))
    \_al_u2040|_al_u2127  (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_6 ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/n576 [28],\picorv32_core/n576 [20]}),
    .c({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_prefetch_placeOpt_6 }),
    .d({_al_u1546_o_placeOpt_3,_al_u1546_o_placeOpt_3}),
    .f({_al_u2040_o,_al_u2127_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTF1("~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("(B*~(~1*~(~A*~(C*~D))))"),
    //.LUTG1("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0100010000000100),
    .INIT_LUTF1(16'b0101010001010100),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b0101000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2042|_al_u2041  (
    .a({\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_4 ,\picorv32_core/n669_lutinv_placeOpt_3 }),
    .c({\picorv32_core/mem_do_wdata ,\picorv32_core/mem_do_prefetch_placeOpt_4 }),
    .d({open_n12264,_al_u1546_o_placeOpt_5}),
    .e({_al_u1546_o_placeOpt_5,\picorv32_core/pcpi_rs1$28$ }),
    .f({_al_u2042_o,_al_u2041_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(A*~(~1*~B*~(C*~D)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2043 (
    .a({\picorv32_core/n668_lutinv ,\picorv32_core/mem_do_prefetch_placeOpt_4 }),
    .b({\picorv32_core/n576 [28],\picorv32_core/n576 [28]}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_4 ,\picorv32_core/n668_lutinv }),
    .d({_al_u1546_o_placeOpt_5,_al_u1546_o_placeOpt_5}),
    .mi({open_n12297,\picorv32_core/mem_do_wdata }),
    .fx({open_n12302,_al_u2043_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*A*~(B*~(0*~D)))"),
    //.LUT1("(~C*A*~(B*~(1*~D)))"),
    .INIT_LUT0(16'b0000001000000010),
    .INIT_LUT1(16'b0000001000001010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2045 (
    .a({\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv ,\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv }),
    .b({_al_u2014_o,_al_u2014_o}),
    .c({_al_u2044_o,_al_u2044_o}),
    .d({_al_u1302_o,_al_u1302_o}),
    .mi({open_n12317,\picorv32_core/pcpi_rs1$24$ }),
    .fx({open_n12322,_al_u2045_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~D*B*C*~A+~D*B*C*A"),
    //.LUTG0("A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG1("D*B*~C*~A+~D*B*C*~A+D*B*C*~A+D*B*~C*A+~D*B*C*A+D*B*C*A"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b1010101000000000),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2046|_al_u2142  (
    .a({open_n12325,\picorv32_core/cpuregs_p1/dram_do_i1_001 }),
    .b({_al_u1926_o,open_n12326}),
    .c({\picorv32_core/cpuregs_p1/dram_do_i0_028 ,\picorv32_core/cpuregs_p1/dram_do_i0_001 }),
    .d({\picorv32_core/decoded_rs1 [4],_al_u1926_o}),
    .e({\picorv32_core/cpuregs_p1/dram_do_i1_028 ,\picorv32_core/decoded_rs1 [4]}),
    .f({_al_u2046_o,_al_u2142_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("(~D*~A*~B*~(0*~C))"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("(~D*~A*~B*~(1*~C))"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0000000000010001),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0000000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2048|_al_u2047  (
    .a({\picorv32_core/sel41_b28/B5 ,_al_u2046_o}),
    .b({_al_u2045_o,\picorv32_core/n664_lutinv_placeOpt_7 }),
    .c({_al_u1924_o,\picorv32_core/instr_lui }),
    .d({\picorv32_core/sel43_b28/B2 ,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/reg_pc [28]}),
    .f({_al_u2048_o,\picorv32_core/sel41_b28/B5 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~B*~C*~A*~D+B*~C*~A*~D+~B*~C*~A*D+B*~C*~A*D+~B*~C*A*D+B*~C*A*D"),
    //.LUTG0("0"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0101010100000101),
    .INIT_LUTF1(16'b0000111100000101),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2050|_al_u2094  (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_7 ,\picorv32_core/mem_do_rdata }),
    .c({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .d({_al_u1546_o_placeOpt_7,_al_u1546_o_placeOpt_7}),
    .e({\picorv32_core/n576 [27],\picorv32_core/n576 [23]}),
    .f({_al_u2050_o,_al_u2094_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUT1("(B*~(~1*~(~A*~(C*~D))))"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b1100110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2051 (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/n669_lutinv_placeOpt_4 ,\picorv32_core/n669_lutinv_placeOpt_4 }),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_7 ,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .d({_al_u1546_o_placeOpt_1,_al_u1546_o_placeOpt_1}),
    .mi({open_n12407,\picorv32_core/pcpi_rs1$27$ }),
    .fx({open_n12412,_al_u2051_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(A*~(~1*~B*~(D*~C)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2053 (
    .a({\picorv32_core/n668_lutinv ,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .b({\picorv32_core/n576 [27],\picorv32_core/n576 [27]}),
    .c({_al_u1546_o_placeOpt_1,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/mem_do_prefetch_placeOpt_7 ,_al_u1546_o_placeOpt_1}),
    .mi({open_n12427,\picorv32_core/mem_do_wdata }),
    .fx({open_n12432,_al_u2053_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010110000000000),
    .MODE("LOGIC"))
    \_al_u2054|_al_u2131  (
    .a({\picorv32_core/cpuregs_p1/dram_do_i1_027 ,_al_u1926_o}),
    .b({\picorv32_core/cpuregs_p1/dram_do_i0_027 ,\picorv32_core/decoded_rs1 [4]}),
    .c({\picorv32_core/decoded_rs1 [4],\picorv32_core/cpuregs_p1/dram_do_i0_020 }),
    .d({_al_u1926_o,\picorv32_core/cpuregs_p1/dram_do_i1_020 }),
    .f({_al_u2054_o,_al_u2131_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(C*~(~A*~(1*B*~D)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010000011100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2055 (
    .a({_al_u2054_o,_al_u2054_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv_placeOpt_3 }),
    .c({\picorv32_core/n664_lutinv_placeOpt_3 ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/instr_lui ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n12467,\picorv32_core/reg_pc [27]}),
    .fx({open_n12472,\picorv32_core/sel41_b27/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*~(B*~D)))"),
    //.LUT1("(~A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUT0(16'b0101000001010100),
    .INIT_LUT1(16'b0001000100000101),
    .MODE("LOGIC"))
    \_al_u2056|_al_u2063  (
    .a({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$26$ }),
    .b({\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/mem_do_prefetch_placeOpt_3 }),
    .c({\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/mem_do_wdata }),
    .d({_al_u1302_o,_al_u1546_o_placeOpt_4}),
    .f({_al_u2056_o,_al_u2063_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b0010001000001010),
    .MODE("LOGIC"))
    \_al_u2057|_al_u2089  (
    .a({\picorv32_core/n554 ,\picorv32_core/n554 }),
    .b({\picorv32_core/pcpi_rs1$31$ ,_al_u1302_o}),
    .c({\picorv32_core/pcpi_rs1$23$ ,\picorv32_core/pcpi_rs1$23$ }),
    .d({_al_u1302_o,\picorv32_core/pcpi_rs1$25$ }),
    .f({_al_u2057_o,_al_u2089_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUTF1("(~D*~B*~(A*~C))"),
    //.LUTG0("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    //.LUTG1("(~D*~B*~(A*~C))"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000110001),
    .INIT_LUTG0(16'b1010101000000010),
    .INIT_LUTG1(16'b0000000000110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2059|_al_u2058  (
    .a({\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/n667_lutinv }),
    .b({\picorv32_core/sel41_b27/B5 ,_al_u2056_o}),
    .c({_al_u1924_o,_al_u2057_o}),
    .d({\picorv32_core/sel41_b27/B2 ,_al_u1313_o}),
    .e({open_n12517,\picorv32_core/pcpi_rs1$27$ }),
    .f({_al_u2059_o,\picorv32_core/sel41_b27/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~D*~A*~C*~B+~D*A*~C*~B+~D*~A*C*~B+~D*A*C*~B+~D*~A*C*B+~D*A*C*B"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2061|_al_u2064  (
    .a({open_n12538,\picorv32_core/mem_do_prefetch_placeOpt_3 }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_3 ,\picorv32_core/n576 [26]}),
    .c({_al_u1546_o_placeOpt_3,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/mem_do_rdata ,_al_u1546_o_placeOpt_3}),
    .e({\picorv32_core/n576 [26],\picorv32_core/mem_do_wdata }),
    .f({_al_u2061_o,_al_u2064_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUT1("(A*~(~1*~(~C*~(B*~D))))"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2062 (
    .a({\picorv32_core/n669_lutinv_placeOpt_3 ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_3 ,\picorv32_core/n669_lutinv_placeOpt_3 }),
    .c({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_prefetch_placeOpt_3 }),
    .d({_al_u1546_o_placeOpt_4,_al_u1546_o_placeOpt_4}),
    .mi({open_n12573,\picorv32_core/pcpi_rs1$26$ }),
    .fx({open_n12578,_al_u2062_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1100000010100000),
    .MODE("LOGIC"))
    \_al_u2065|_al_u2120  (
    .a({\picorv32_core/cpuregs_p1/dram_do_i0_026 ,_al_u1926_o}),
    .b({\picorv32_core/cpuregs_p1/dram_do_i1_026 ,\picorv32_core/decoded_rs1 [4]}),
    .c({_al_u1926_o,\picorv32_core/cpuregs_p1/dram_do_i0_021 }),
    .d({\picorv32_core/decoded_rs1 [4],\picorv32_core/cpuregs_p1/dram_do_i1_021 }),
    .f({_al_u2065_o,_al_u2120_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(C*~(~A*~(1*B*~D)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010000011100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2066 (
    .a({_al_u2065_o,_al_u2065_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv_placeOpt_3 }),
    .c({\picorv32_core/n664_lutinv_placeOpt_3 ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/instr_lui ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n12613,\picorv32_core/reg_pc [26]}),
    .fx({open_n12618,\picorv32_core/sel41_b26/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*~(B*~D)))"),
    //.LUT1("(~A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUT0(16'b0101000001010100),
    .INIT_LUT1(16'b0001000100000101),
    .MODE("LOGIC"))
    \_al_u2067|_al_u2074  (
    .a({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$25$ }),
    .b({\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/mem_do_prefetch_placeOpt_4 }),
    .c({\picorv32_core/pcpi_rs1$25$ ,\picorv32_core/mem_do_wdata }),
    .d({_al_u1302_o,_al_u1546_o_placeOpt_3}),
    .f({_al_u2067_o,_al_u2074_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b0010001000001010),
    .MODE("LOGIC"))
    \_al_u2068|_al_u2100  (
    .a({\picorv32_core/n554 ,\picorv32_core/n554 }),
    .b({\picorv32_core/pcpi_rs1$30$ ,_al_u1302_o}),
    .c({\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs1$22$ }),
    .d({_al_u1302_o,\picorv32_core/pcpi_rs1$24$ }),
    .f({_al_u2068_o,_al_u2100_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    //.LUTG0("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b1010101000000010),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2070|_al_u2069  (
    .a({open_n12661,\picorv32_core/n667_lutinv }),
    .b({\picorv32_core/sel41_b26/B5 ,_al_u2067_o}),
    .c({_al_u1924_o,_al_u2068_o}),
    .d({\picorv32_core/sel41_b26/B2 ,_al_u1313_o}),
    .e({\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$26$ }),
    .f({_al_u2070_o,\picorv32_core/sel41_b26/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~A*~C*~B*~D+~A*~C*B*~D"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*~C*B*~D+A*~C*B*~D"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000000000101),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2072|_al_u2075  (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_4 ,\picorv32_core/mem_do_prefetch_placeOpt_4 }),
    .b({open_n12684,\picorv32_core/n576 [25]}),
    .c({\picorv32_core/n576 [25],\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/mem_do_rdata ,_al_u1546_o_placeOpt_5}),
    .e({_al_u1546_o_placeOpt_5,\picorv32_core/mem_do_wdata }),
    .f({_al_u2072_o,_al_u2075_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(A*~C)*~(D*~B))"),
    //.LUTF1("(A*~(~0*~(~D*~(B*~C))))"),
    //.LUTG0("~(1*~(A*~C)*~(D*~B))"),
    //.LUTG1("(A*~(~1*~(~D*~(B*~C))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0000000010100010),
    .INIT_LUTG0(16'b0011101100001010),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2073|picorv32_core/reg25_b25  (
    .a({\picorv32_core/n669_lutinv_placeOpt_3 ,_al_u2075_o}),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_4 ,_al_u2072_o}),
    .c({_al_u1546_o_placeOpt_3,_al_u2074_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_do_rdata ,_al_u2073_o}),
    .e({\picorv32_core/pcpi_rs1$25$ ,_al_u2081_o}),
    .f({_al_u2073_o,open_n12722}),
    .q({open_n12726,\picorv32_core/pcpi_rs1$25$ }));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("0"),
    //.LUTG0("~C*~B*A*~D+C*~B*A*~D+~C*B*~A*D+C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG1("~D*~B*A*~C+D*~B*A*~C+~D*B*~A*C+D*B*~A*C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1110111000100010),
    .INIT_LUTG1(16'b1110001011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2076|_al_u2109  (
    .a({\picorv32_core/cpuregs_p1/dram_do_i0_025 ,\picorv32_core/cpuregs_p1/dram_do_i0_022 }),
    .b({\picorv32_core/decoded_rs1 [4],\picorv32_core/decoded_rs1 [4]}),
    .c({\picorv32_core/cpuregs_p1/dram_do_i1_025 ,open_n12727}),
    .d({open_n12730,\picorv32_core/cpuregs_p1/dram_do_i1_022 }),
    .e({_al_u1926_o,_al_u1926_o}),
    .f({_al_u2076_o,_al_u2109_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*B*~A*~C+~D*~B*A*~C+~D*B*A*~C+~D*B*~A*C+~D*~B*A*C+~D*B*A*C"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D"),
    //.LUTG0("~D*~B*A*~C+~D*B*A*~C+~D*~B*A*C+~D*B*A*C"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000011101110),
    .INIT_LUTF1(16'b0000010110101111),
    .INIT_LUTG0(16'b0000000010101010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2078|_al_u2085  (
    .a({_al_u1302_o,\picorv32_core/mem_do_wdata }),
    .b({open_n12751,\picorv32_core/mem_do_prefetch_placeOpt_4 }),
    .c({\picorv32_core/pcpi_rs1$24$ ,open_n12752}),
    .d({\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$24$ }),
    .e({\picorv32_core/n554 ,_al_u1546_o_placeOpt_5}),
    .f({_al_u2078_o,_al_u2085_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~D*~C+~A*~B*D*~C+~A*B*D*~C+~A*B*~D*C+~A*~B*D*C+~A*B*D*C"),
    //.LUTF1("A*~B*~D*~C+A*~B*D*~C+A*B*D*~C+A*~B*~D*C+A*~B*D*C+A*B*D*C"),
    //.LUTG0("~A*~B*D*~C+~A*B*D*~C+~A*~B*D*C+~A*B*D*C"),
    //.LUTG1("A*~B*~D*~C+A*~B*~D*C"),
    .INIT_LUTF0(16'b0101010101000100),
    .INIT_LUTF1(16'b1010101000100010),
    .INIT_LUTG0(16'b0101010100000000),
    .INIT_LUTG1(16'b0000000000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2079|_al_u2118  (
    .a({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$21$ }),
    .b({\picorv32_core/pcpi_rs1$21$ ,\picorv32_core/mem_do_prefetch_placeOpt_3 }),
    .d({_al_u1302_o,\picorv32_core/mem_do_wdata }),
    .e({\picorv32_core/pcpi_rs1$29$ ,_al_u1546_o_placeOpt_4}),
    .f({_al_u2079_o,_al_u2118_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUT1("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2080 (
    .a({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .b({_al_u2078_o,_al_u2078_o}),
    .c({_al_u2079_o,_al_u2079_o}),
    .d({_al_u1313_o,_al_u1313_o}),
    .mi({open_n12811,\picorv32_core/pcpi_rs1$25$ }),
    .fx({open_n12816,\picorv32_core/sel41_b25/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("~A*~B*~D*~C+~A*~B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("~A*~B*D*~C+~A*~B*D*C"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0001000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2081|_al_u2077  (
    .a({\picorv32_core/sel41_b25/B5 ,_al_u2076_o}),
    .b({\picorv32_core/sel41_b25/B2 ,\picorv32_core/n664_lutinv_placeOpt_3 }),
    .c({open_n12819,\picorv32_core/instr_lui }),
    .d({_al_u1924_o,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/pcpi_rs1$25$ ,\picorv32_core/reg_pc [25]}),
    .f({_al_u2081_o,\picorv32_core/sel41_b25/B5 }));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(D*~B)*~(A*~C))"),
    //.LUTF1("(A*~(~0*~(~D*~(B*~C))))"),
    //.LUTG0("~(1*~(D*~B)*~(A*~C))"),
    //.LUTG1("(A*~(~1*~(~D*~(B*~C))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0000000010100010),
    .INIT_LUTG0(16'b0011101100001010),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2084|picorv32_core/reg25_b24  (
    .a({\picorv32_core/n669_lutinv_placeOpt_3 ,_al_u2084_o}),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_4 ,_al_u2085_o}),
    .c({_al_u1546_o_placeOpt_5,_al_u2083_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_do_rdata ,_al_u2086_o}),
    .e({\picorv32_core/pcpi_rs1$24$ ,_al_u2092_o}),
    .f({_al_u2084_o,open_n12857}),
    .q({open_n12861,\picorv32_core/pcpi_rs1$24$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(C*~(~1*~B*~(A*~D)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2086 (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_4 ,\picorv32_core/mem_do_prefetch_placeOpt_4 }),
    .b({\picorv32_core/n576 [24],\picorv32_core/n576 [24]}),
    .c({\picorv32_core/n668_lutinv ,\picorv32_core/n668_lutinv }),
    .d({_al_u1546_o_placeOpt_5,_al_u1546_o_placeOpt_5}),
    .mi({open_n12874,\picorv32_core/mem_do_wdata }),
    .fx({open_n12879,_al_u2086_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*C*~D+A*B*C*~D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("A*B*~C*D+A*B*C*D"),
    //.LUTG0("A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG1("A*~B*~C*~D+A*~B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1010000010100000),
    .INIT_LUTF1(16'b1000100000000000),
    .INIT_LUTG0(16'b1010101000000000),
    .INIT_LUTG1(16'b1010101000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2087|_al_u2098  (
    .a({_al_u1926_o,_al_u1926_o}),
    .b({\picorv32_core/decoded_rs1 [4],open_n12882}),
    .c({open_n12883,\picorv32_core/cpuregs_p1/dram_do_i0_023 }),
    .d({\picorv32_core/cpuregs_p1/dram_do_i1_024 ,\picorv32_core/cpuregs_p1/dram_do_i1_023 }),
    .e({\picorv32_core/cpuregs_p1/dram_do_i0_024 ,\picorv32_core/decoded_rs1 [4]}),
    .f({_al_u2087_o,_al_u2098_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*~(B*~D)))"),
    //.LUT1("(A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUT0(16'b0101000001010100),
    .INIT_LUT1(16'b0010001000001010),
    .MODE("LOGIC"))
    \_al_u2090|_al_u2129  (
    .a({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$20$ }),
    .b({\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/mem_do_prefetch_placeOpt_3 }),
    .c({\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/mem_do_wdata }),
    .d({_al_u1302_o,_al_u1546_o_placeOpt_3}),
    .f({_al_u2090_o,_al_u2129_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUT1("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2091 (
    .a({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .b({_al_u2089_o,_al_u2089_o}),
    .c({_al_u2090_o,_al_u2090_o}),
    .d({_al_u1313_o,_al_u1313_o}),
    .mi({open_n12938,\picorv32_core/pcpi_rs1$24$ }),
    .fx({open_n12943,\picorv32_core/sel41_b24/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0000000000000101),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2092|_al_u2088  (
    .a({\picorv32_core/pcpi_rs1$24$ ,_al_u2087_o}),
    .b({open_n12946,\picorv32_core/n664_lutinv_placeOpt_3 }),
    .c({\picorv32_core/sel41_b24/B2 ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/sel41_b24/B5 ,\picorv32_core/is_lui_auipc_jal }),
    .e({_al_u1924_o,\picorv32_core/reg_pc [24]}),
    .f({_al_u2092_o,\picorv32_core/sel41_b24/B5 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTF1("~D*B*~A*~C+~D*~B*A*~C+~D*B*A*~C+~D*B*~A*C+~D*~B*A*C+~D*B*A*C"),
    //.LUTG0("(B*~(~1*~(~A*~(C*~D))))"),
    //.LUTG1("~D*~B*A*~C+~D*B*A*~C+~D*~B*A*C+~D*B*A*C"),
    .INIT_LUTF0(16'b0100010000000100),
    .INIT_LUTF1(16'b0000000011101110),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b0000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2096|_al_u2095  (
    .a({\picorv32_core/mem_do_wdata ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_7 ,\picorv32_core/n669_lutinv_placeOpt_2 }),
    .c({open_n12969,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .d({\picorv32_core/pcpi_rs1$23$ ,_al_u1546_o_placeOpt_7}),
    .e({_al_u1546_o_placeOpt_7,\picorv32_core/pcpi_rs1$23$ }),
    .f({_al_u2096_o,_al_u2095_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(A*~(~1*~D*~(B*~C)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2097 (
    .a({\picorv32_core/n668_lutinv ,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_7 ,\picorv32_core/n576 [23]}),
    .c({_al_u1546_o_placeOpt_7,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/n576 [23],_al_u1546_o_placeOpt_7}),
    .mi({open_n13004,\picorv32_core/mem_do_wdata }),
    .fx({open_n13009,_al_u2097_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(D*~(~A*~(1*B*~C)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010111000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2099 (
    .a({_al_u2098_o,_al_u2098_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv_placeOpt_3 }),
    .c({\picorv32_core/instr_lui ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/n664_lutinv_placeOpt_3 ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n13024,\picorv32_core/reg_pc [23]}),
    .fx({open_n13029,\picorv32_core/sel41_b23/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*~(B*~D)))"),
    //.LUT1("(A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUT0(16'b0101000001010100),
    .INIT_LUT1(16'b0000001010001010),
    .MODE("LOGIC"))
    \_al_u2101|_al_u2150  (
    .a({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$19$ }),
    .b({_al_u1302_o,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .c({\picorv32_core/pcpi_rs1$19$ ,\picorv32_core/mem_do_wdata }),
    .d({\picorv32_core/pcpi_rs1$27$ ,_al_u1546_o_placeOpt_2}),
    .f({_al_u2101_o,_al_u2150_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUTF1("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG0("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0100010001010101),
    .INIT_LUTG0(16'b1010101000000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2103|_al_u2102  (
    .a({\picorv32_core/sel41_b23/B2 ,\picorv32_core/n667_lutinv }),
    .b({_al_u1924_o,_al_u2100_o}),
    .c({open_n13052,_al_u2101_o}),
    .d({\picorv32_core/pcpi_rs1$23$ ,_al_u1313_o}),
    .e({\picorv32_core/sel41_b23/B5 ,\picorv32_core/pcpi_rs1$23$ }),
    .f({_al_u2103_o,\picorv32_core/sel41_b23/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~C*~D*~B*~A+~C*~D*~B*A"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~C*~D*~B*~A+~C*~D*B*~A+~C*~D*~B*A+~C*~D*B*A"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2105|_al_u2108  (
    .a({open_n13075,\picorv32_core/mem_do_prefetch_placeOpt_3 }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_3 ,\picorv32_core/n576 [22]}),
    .c({\picorv32_core/mem_do_rdata ,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/n576 [22],_al_u1546_o_placeOpt_4}),
    .e({_al_u1546_o_placeOpt_4,\picorv32_core/mem_do_wdata }),
    .f({_al_u2105_o,_al_u2108_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTF1("~D*B*~A*~C+~D*~B*A*~C+~D*B*A*~C+~D*B*~A*C+~D*~B*A*C+~D*B*A*C"),
    //.LUTG0("(B*~(~1*~(~A*~(C*~D))))"),
    //.LUTG1("~D*~B*A*~C+~D*B*A*~C+~D*~B*A*C+~D*B*A*C"),
    .INIT_LUTF0(16'b0100010000000100),
    .INIT_LUTF1(16'b0000000011101110),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b0000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2107|_al_u2106  (
    .a({\picorv32_core/mem_do_wdata ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/n669_lutinv_placeOpt_2 }),
    .c({open_n13098,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .d({\picorv32_core/pcpi_rs1$22$ ,_al_u1546_o_placeOpt_2}),
    .e({_al_u1546_o_placeOpt_2,\picorv32_core/pcpi_rs1$22$ }),
    .f({_al_u2107_o,_al_u2106_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(C*~(~A*~(1*B*~D)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010000011100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2110 (
    .a({_al_u2109_o,_al_u2109_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv_placeOpt_4 }),
    .c({\picorv32_core/n664_lutinv_placeOpt_4 ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/instr_lui ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n13133,\picorv32_core/reg_pc [22]}),
    .fx({open_n13138,\picorv32_core/sel41_b22/B5 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D"),
    //.LUTF1("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG0("0"),
    //.LUTG1("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT_LUTF0(16'b0000001111001111),
    .INIT_LUTF1(16'b0000000100110001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2111|_al_u2133  (
    .a({\picorv32_core/pcpi_rs1$21$ ,open_n13141}),
    .b({\picorv32_core/n554 ,_al_u1302_o}),
    .c({_al_u1302_o,\picorv32_core/pcpi_rs1$19$ }),
    .d({\picorv32_core/pcpi_rs1$23$ ,\picorv32_core/pcpi_rs1$21$ }),
    .e({open_n13144,\picorv32_core/n554 }),
    .f({_al_u2111_o,_al_u2133_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*B*~A*~C+~D*~B*A*~C+~D*B*A*~C+~D*B*~A*C+~D*~B*A*C+~D*B*A*C"),
    //.LUTF1("D*~B*~C*~A+D*B*~C*~A+D*B*C*~A+D*~B*~C*A+D*B*~C*A+D*B*C*A"),
    //.LUTG0("~D*~B*A*~C+~D*B*A*~C+~D*~B*A*C+~D*B*A*C"),
    //.LUTG1("D*~B*~C*~A+D*~B*~C*A"),
    .INIT_LUTF0(16'b0000000011101110),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b0000000010101010),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2112|_al_u2161  (
    .a({open_n13165,\picorv32_core/mem_do_wdata }),
    .b({_al_u1302_o,\picorv32_core/mem_do_prefetch_placeOpt_3 }),
    .c({\picorv32_core/pcpi_rs1$18$ ,open_n13166}),
    .d({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$18$ }),
    .e({\picorv32_core/pcpi_rs1$26$ ,_al_u1546_o_placeOpt_4}),
    .f({_al_u2112_o,_al_u2161_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUTF1("~A*~B*~C*~D+~A*~B*C*~D"),
    //.LUTG0("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    //.LUTG1("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000010001),
    .INIT_LUTG0(16'b1010101000000010),
    .INIT_LUTG1(16'b0001000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2114|_al_u2113  (
    .a({\picorv32_core/sel41_b22/B2 ,\picorv32_core/n667_lutinv }),
    .b({\picorv32_core/sel41_b22/B5 ,_al_u2111_o}),
    .c({open_n13189,_al_u2112_o}),
    .d({\picorv32_core/pcpi_rs1$22$ ,_al_u1313_o}),
    .e({_al_u1924_o,\picorv32_core/pcpi_rs1$22$ }),
    .f({_al_u2114_o,\picorv32_core/sel41_b22/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~B*~C*~A*~D+~B*C*~A*~D+~B*~C*~A*D+B*~C*~A*D+~B*C*~A*D+B*C*~A*D"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0101010100010001),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2116|_al_u2119  (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_prefetch_placeOpt_3 }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_3 ,\picorv32_core/n576 [21]}),
    .c({open_n13212,\picorv32_core/n668_lutinv }),
    .d({_al_u1546_o_placeOpt_6,_al_u1546_o_placeOpt_6}),
    .e({\picorv32_core/n576 [21],\picorv32_core/mem_do_wdata }),
    .f({_al_u2116_o,_al_u2119_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(D*~A)*~(B*~C))"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~(1*~(D*~A)*~(B*~C))"),
    //.LUTG1("A*B*~C*~D+A*B*C*~D+A*B*~C*D+A*B*C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b1100100011001100),
    .INIT_LUTG0(16'b0101110100001100),
    .INIT_LUTG1(16'b1000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2117|picorv32_core/reg25_b21  (
    .a({\picorv32_core/pcpi_rs1$21$ ,_al_u2118_o}),
    .b({\picorv32_core/n669_lutinv_placeOpt_3 ,_al_u2117_o}),
    .c({_al_u1546_o_placeOpt_4,_al_u2116_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_do_prefetch_placeOpt_3 ,_al_u2119_o}),
    .e({\picorv32_core/mem_do_rdata ,_al_u2125_o}),
    .f({_al_u2117_o,open_n13250}),
    .q({open_n13254,\picorv32_core/pcpi_rs1$21$ }));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~D*~C+~A*B*~D*~C+~A*~B*D*~C+~A*B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    //.LUTF1("~A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D"),
    //.LUTG0("~A*B*~D*~C+~A*B*D*~C"),
    //.LUTG1("~A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D"),
    .INIT_LUTF0(16'b0001010100010101),
    .INIT_LUTF1(16'b0000000100110001),
    .INIT_LUTG0(16'b0000010000000100),
    .INIT_LUTG1(16'b0000000100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2122|_al_u2154  (
    .a({\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/n554 }),
    .b({\picorv32_core/n554 ,_al_u1302_o}),
    .c({_al_u1302_o,\picorv32_core/pcpi_rs1$20$ }),
    .d({\picorv32_core/pcpi_rs1$22$ ,open_n13257}),
    .e({open_n13258,\picorv32_core/pcpi_rs1$18$ }),
    .f({_al_u2122_o,_al_u2154_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*B*~A*~D+C*B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("~A*C*~D*~B+A*C*~D*~B+A*C*D*~B+~A*C*~D*B+A*C*~D*B+A*C*D*B"),
    //.LUTG0("0"),
    //.LUTG1("~A*C*~D*~B+~A*C*~D*B"),
    .INIT_LUTF0(16'b1010101011101110),
    .INIT_LUTF1(16'b1010000011110000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2123|_al_u2172  (
    .a({_al_u1302_o,\picorv32_core/mem_do_wdata }),
    .b({open_n13279,\picorv32_core/mem_do_prefetch_placeOpt_3 }),
    .c({\picorv32_core/n554 ,open_n13280}),
    .d({\picorv32_core/pcpi_rs1$17$ ,_al_u1546_o_placeOpt_3}),
    .e({\picorv32_core/pcpi_rs1$25$ ,\picorv32_core/pcpi_rs1$17$ }),
    .f({_al_u2123_o,_al_u2172_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUT1("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2124 (
    .a({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .b({_al_u2122_o,_al_u2122_o}),
    .c({_al_u2123_o,_al_u2123_o}),
    .d({_al_u1313_o,_al_u1313_o}),
    .mi({open_n13315,\picorv32_core/pcpi_rs1$21$ }),
    .fx({open_n13320,\picorv32_core/sel41_b21/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("~A*~B*~D*~C+~A*~B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("~A*~B*D*~C+~A*~B*D*C"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0001000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2125|_al_u2121  (
    .a({\picorv32_core/sel41_b21/B5 ,_al_u2120_o}),
    .b({\picorv32_core/sel41_b21/B2 ,\picorv32_core/n664_lutinv_placeOpt_4 }),
    .c({open_n13323,\picorv32_core/instr_lui }),
    .d({_al_u1924_o,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/pcpi_rs1$21$ ,\picorv32_core/reg_pc [21]}),
    .f({_al_u2125_o,\picorv32_core/sel41_b21/B5 }));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(D*~C)*~(A*~B))"),
    //.LUTF1("(A*~(~0*~(~D*~(B*~C))))"),
    //.LUTG0("~(1*~(D*~C)*~(A*~B))"),
    //.LUTG1("(A*~(~1*~(~D*~(B*~C))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0000000010100010),
    .INIT_LUTG0(16'b0010111100100010),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2128|picorv32_core/reg25_b20  (
    .a({\picorv32_core/n669_lutinv_placeOpt_3 ,_al_u2128_o}),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_6 ,_al_u2127_o}),
    .c({_al_u1546_o_placeOpt_3,_al_u2129_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_do_rdata ,_al_u2130_o}),
    .e({\picorv32_core/pcpi_rs1$20$ ,_al_u2136_o}),
    .f({_al_u2128_o,open_n13361}),
    .q({open_n13365,\picorv32_core/pcpi_rs1$20$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(B*~(~1*~A*~(C*~D)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1100110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2130 (
    .a({\picorv32_core/n576 [20],\picorv32_core/mem_do_prefetch_placeOpt_6 }),
    .b({\picorv32_core/n668_lutinv ,\picorv32_core/n576 [20]}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_6 ,\picorv32_core/n668_lutinv }),
    .d({_al_u1546_o_placeOpt_3,_al_u1546_o_placeOpt_3}),
    .mi({open_n13378,\picorv32_core/mem_do_wdata }),
    .fx({open_n13383,_al_u2130_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b0000001010100010),
    .MODE("LOGIC"))
    \_al_u2134|_al_u2176  (
    .a({\picorv32_core/n554 ,\picorv32_core/n554 }),
    .b({\picorv32_core/pcpi_rs1$16$ ,_al_u1302_o}),
    .c({_al_u1302_o,\picorv32_core/pcpi_rs1$16$ }),
    .d({\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/pcpi_rs1$18$ }),
    .f({_al_u2134_o,_al_u2176_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUT1("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2135 (
    .a({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .b({_al_u2133_o,_al_u2133_o}),
    .c({_al_u2134_o,_al_u2134_o}),
    .d({_al_u1313_o,_al_u1313_o}),
    .mi({open_n13418,\picorv32_core/pcpi_rs1$20$ }),
    .fx({open_n13423,\picorv32_core/sel41_b20/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0000000000001101),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0000000000001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2136|_al_u2132  (
    .a({\picorv32_core/pcpi_rs1$20$ ,_al_u2131_o}),
    .b({_al_u1924_o,\picorv32_core/n664_lutinv_placeOpt_4 }),
    .c({\picorv32_core/sel41_b20/B2 ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/sel41_b20/B5 ,\picorv32_core/is_lui_auipc_jal }),
    .e({open_n13428,\picorv32_core/reg_pc [20]}),
    .f({_al_u2136_o,\picorv32_core/sel41_b20/B5 }));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(C*~B)*~(A*~D))"),
    //.LUTF1("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTG0("~(1*~(C*~B)*~(A*~D))"),
    //.LUTG1("(B*~(~1*~(~A*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0100010000000100),
    .INIT_LUTG0(16'b0011000010111010),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2139|picorv32_core/reg25_b1  (
    .a({\picorv32_core/mem_do_rdata ,_al_u2139_o}),
    .b({\picorv32_core/n669_lutinv_placeOpt_2 ,_al_u2140_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_7 ,_al_u2141_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o_placeOpt_1,_al_u2138_o}),
    .e({\picorv32_core/pcpi_rs1$1$ ,_al_u2146_o}),
    .f({_al_u2139_o,open_n13464}),
    .q({open_n13468,\picorv32_core/pcpi_rs1$1$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~0*~C*~(A*~D)))"),
    //.LUT1("(B*~(~1*~C*~(A*~D)))"),
    .INIT_LUT0(16'b1100000011001000),
    .INIT_LUT1(16'b1100110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2141 (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_7 ,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .b({\picorv32_core/n668_lutinv ,\picorv32_core/n668_lutinv }),
    .c({\picorv32_core/n576 [1],\picorv32_core/n576 [1]}),
    .d({_al_u1546_o_placeOpt_1,_al_u1546_o_placeOpt_1}),
    .mi({open_n13481,\picorv32_core/mem_do_wdata }),
    .fx({open_n13486,_al_u2141_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~D*~(0*A*~C)))"),
    //.LUT1("(A*~(~D*~(1*B*~C)))"),
    .INIT_LUT0(16'b1100110000000000),
    .INIT_LUT1(16'b1010101000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2143 (
    .a({\picorv32_core/n664_lutinv_placeOpt_7 ,\picorv32_core/is_lui_auipc_jal }),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv_placeOpt_7 }),
    .c({\picorv32_core/instr_lui ,\picorv32_core/instr_lui }),
    .d({_al_u2142_o,_al_u2142_o}),
    .mi({open_n13501,\picorv32_core/reg_pc [1]}),
    .fx({open_n13506,\picorv32_core/sel41_b1/B5 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+~(A)*B*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+A*B*~(C)*D*~(0)+A*~(B)*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("(~C*~(B*(~A*~(0)*~(D)+~A*0*~(D)+~(~A)*0*D+~A*0*D)))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+~(A)*B*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+A*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+A*B*~(C)*D*~(1)+A*~(B)*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("(~C*~(B*(~A*~(1)*~(D)+~A*1*~(D)+~(~A)*1*D+~A*1*D)))"),
    .INIT_LUTF0(16'b1010101111101111),
    .INIT_LUTF1(16'b0000111100001011),
    .INIT_LUTG0(16'b0010001101100111),
    .INIT_LUTG1(16'b0000001100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2145|_al_u2144  (
    .a({_al_u2144_o,\picorv32_core/n554 }),
    .b({\picorv32_core/n667_lutinv ,_al_u1302_o}),
    .c({\picorv32_core/sel41_b1/B5 ,\picorv32_core/pcpi_rs1$0$ }),
    .d({_al_u1313_o,\picorv32_core/pcpi_rs1$2$ }),
    .e({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$5$ }),
    .f({_al_u2145_o,_al_u2144_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTF1("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0101000001010000),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1111000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2146|_al_u1997  (
    .a({\picorv32_core/pcpi_rs1$1$ ,open_n13531}),
    .c({_al_u2145_o,\picorv32_core/pcpi_rs1$3$ }),
    .d({open_n13536,_al_u1996_o}),
    .e({_al_u1924_o,_al_u1924_o}),
    .f({_al_u2146_o,_al_u1997_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~A*~D*~C*~B+~A*~D*~C*B"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~A*~D*~C*~B+~A*~D*C*~B+~A*~D*~C*B+~A*~D*C*B"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000000000101),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2148|_al_u2151  (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .b({open_n13557,\picorv32_core/n576 [19]}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/n576 [19],_al_u1546_o_placeOpt_2}),
    .e({_al_u1546_o_placeOpt_2,\picorv32_core/mem_do_wdata }),
    .f({_al_u2148_o,_al_u2151_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUT1("(A*~(~1*~(~B*~(C*~D))))"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2149 (
    .a({\picorv32_core/n669_lutinv_placeOpt_2 ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_rdata ,\picorv32_core/n669_lutinv_placeOpt_2 }),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .d({_al_u1546_o_placeOpt_2,_al_u1546_o_placeOpt_2}),
    .mi({open_n13592,\picorv32_core/pcpi_rs1$19$ }),
    .fx({open_n13597,_al_u2149_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(D*~(~A*~(1*B*~C)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010111000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2153 (
    .a({_al_u2152_o,_al_u2152_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv }),
    .c({\picorv32_core/instr_lui ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/n664_lutinv ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n13612,\picorv32_core/reg_pc [19]}),
    .fx({open_n13617,\picorv32_core/sel41_b19/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b0010001000001010),
    .MODE("LOGIC"))
    \_al_u2155|_al_u2187  (
    .a({\picorv32_core/n554 ,\picorv32_core/n554 }),
    .b({\picorv32_core/pcpi_rs1$23$ ,_al_u1302_o}),
    .c({\picorv32_core/pcpi_rs1$15$ ,\picorv32_core/pcpi_rs1$15$ }),
    .d({_al_u1302_o,\picorv32_core/pcpi_rs1$17$ }),
    .f({_al_u2155_o,_al_u2187_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1010101000000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2157|_al_u2156  (
    .a({open_n13640,\picorv32_core/n667_lutinv }),
    .b({\picorv32_core/pcpi_rs1$19$ ,_al_u2154_o}),
    .c({_al_u1924_o,_al_u2155_o}),
    .d({\picorv32_core/sel41_b19/B2 ,_al_u1313_o}),
    .e({\picorv32_core/sel41_b19/B5 ,\picorv32_core/pcpi_rs1$19$ }),
    .f({_al_u2157_o,\picorv32_core/sel41_b19/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~A*~B*~D*~C+~A*~B*D*~C"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~A*~B*~D*~C+~A*~B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000100000001),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0001000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2159|_al_u2162  (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_prefetch_placeOpt_3 }),
    .b({\picorv32_core/n576 [18],\picorv32_core/n576 [18]}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_3 ,\picorv32_core/n668_lutinv }),
    .d({open_n13665,_al_u1546_o_placeOpt_4}),
    .e({_al_u1546_o_placeOpt_4,\picorv32_core/mem_do_wdata }),
    .f({_al_u2159_o,_al_u2162_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUT1("(A*~(~1*~(~C*~(B*~D))))"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2160 (
    .a({\picorv32_core/n669_lutinv_placeOpt_3 ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_3 ,\picorv32_core/n669_lutinv_placeOpt_3 }),
    .c({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_prefetch_placeOpt_3 }),
    .d({_al_u1546_o_placeOpt_4,_al_u1546_o_placeOpt_4}),
    .mi({open_n13698,\picorv32_core/pcpi_rs1$18$ }),
    .fx({open_n13703,_al_u2160_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*((~C*~A)*~(0)*~(D)+(~C*~A)*0*~(D)+~((~C*~A))*0*D+(~C*~A)*0*D))"),
    //.LUTF1("~A*~C*~D*~B+~A*C*~D*~B+~A*~C*~D*B+~A*C*~D*B"),
    //.LUTG0("(B*((~C*~A)*~(1)*~(D)+(~C*~A)*1*~(D)+~((~C*~A))*1*D+(~C*~A)*1*D))"),
    //.LUTG1("~A*~C*~D*~B+~A*~C*D*~B+~A*~C*~D*B+~A*~C*D*B"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b1100110000000100),
    .INIT_LUTG1(16'b0000010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2165|_al_u2167  (
    .a({\picorv32_core/n554 ,_al_u2165_o}),
    .b({open_n13706,\picorv32_core/n667_lutinv }),
    .c({\picorv32_core/pcpi_rs1$19$ ,_al_u2166_o}),
    .d({\picorv32_core/pcpi_rs1$17$ ,_al_u1313_o}),
    .e({_al_u1302_o,\picorv32_core/pcpi_rs1$18$ }),
    .f({_al_u2165_o,\picorv32_core/sel41_b18/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D"),
    //.LUTF1("~C*B*~A*~D+C*B*~A*~D+~C*B*A*~D+C*B*A*~D+~C*B*~A*D+~C*B*A*D"),
    //.LUTG0("A*B*~C*~D+A*B*~C*D"),
    //.LUTG1("C*B*~A*~D+C*B*A*~D"),
    .INIT_LUTF0(16'b0010101000101010),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000100000001000),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2166|_al_u2254  (
    .a({open_n13729,\picorv32_core/n554 }),
    .b({\picorv32_core/n554 ,_al_u1302_o}),
    .c({_al_u1302_o,\picorv32_core/pcpi_rs1$14$ }),
    .d({\picorv32_core/pcpi_rs1$22$ ,open_n13732}),
    .e({\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$6$ }),
    .f({_al_u2166_o,_al_u2254_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0100010001010101),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2168|_al_u2164  (
    .a({\picorv32_core/sel41_b18/B5 ,_al_u2163_o}),
    .b({_al_u1924_o,\picorv32_core/n664_lutinv_placeOpt_2 }),
    .c({open_n13753,\picorv32_core/instr_lui }),
    .d({\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/sel41_b18/B2 ,\picorv32_core/reg_pc [18]}),
    .f({_al_u2168_o,\picorv32_core/sel41_b18/B5 }));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(B*~C)*~(A*~D))"),
    //.LUTF1("(A*~(~0*~(~B*~(C*~D))))"),
    //.LUTG0("~(1*~(B*~C)*~(A*~D))"),
    //.LUTG1("(A*~(~1*~(~B*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0010001000000010),
    .INIT_LUTG0(16'b0000110010101110),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2171|picorv32_core/reg25_b17  (
    .a({\picorv32_core/n669_lutinv_placeOpt_3 ,_al_u2171_o}),
    .b({\picorv32_core/mem_do_rdata ,_al_u2173_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_3 ,_al_u2172_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o_placeOpt_6,_al_u2170_o}),
    .e({\picorv32_core/pcpi_rs1$17$ ,_al_u2179_o}),
    .f({_al_u2171_o,open_n13791}),
    .q({open_n13795,\picorv32_core/pcpi_rs1$17$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(C*~(~1*~B*~(A*~D)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2173 (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_6 ,\picorv32_core/mem_do_prefetch_placeOpt_6 }),
    .b({\picorv32_core/n576 [17],\picorv32_core/n576 [17]}),
    .c({\picorv32_core/n668_lutinv ,\picorv32_core/n668_lutinv }),
    .d({_al_u1546_o_placeOpt_6,_al_u1546_o_placeOpt_6}),
    .mi({open_n13808,\picorv32_core/mem_do_wdata }),
    .fx({open_n13813,_al_u2173_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*~(B*~D)))"),
    //.LUT1("(A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUT0(16'b0101000001010100),
    .INIT_LUT1(16'b0000001010001010),
    .MODE("LOGIC"))
    \_al_u2177|_al_u2216  (
    .a({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$13$ }),
    .b({_al_u1302_o,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .c({\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/mem_do_wdata }),
    .d({\picorv32_core/pcpi_rs1$21$ ,_al_u1546_o_placeOpt_7}),
    .f({_al_u2177_o,_al_u2216_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUT1("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2178 (
    .a({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .b({_al_u2176_o,_al_u2176_o}),
    .c({_al_u2177_o,_al_u2177_o}),
    .d({_al_u1313_o,_al_u1313_o}),
    .mi({open_n13848,\picorv32_core/pcpi_rs1$17$ }),
    .fx({open_n13853,\picorv32_core/sel41_b17/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("~B*~C*~A*~D+B*~C*~A*~D+~B*C*~A*~D+B*C*~A*~D"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("~B*C*~A*~D+B*C*~A*~D"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0000000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2179|_al_u2175  (
    .a({\picorv32_core/sel41_b17/B2 ,_al_u2174_o}),
    .b({open_n13856,\picorv32_core/n664_lutinv_placeOpt_2 }),
    .c({_al_u1924_o,\picorv32_core/instr_lui }),
    .d({\picorv32_core/sel41_b17/B5 ,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/pcpi_rs1$17$ ,\picorv32_core/reg_pc [17]}),
    .f({_al_u2179_o,\picorv32_core/sel41_b17/B5 }));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(C*~B)*~(A*~D))"),
    //.LUTF1("(A*~(~0*~(~B*~(C*~D))))"),
    //.LUTG0("~(1*~(C*~B)*~(A*~D))"),
    //.LUTG1("(A*~(~1*~(~B*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0010001000000010),
    .INIT_LUTG0(16'b0011000010111010),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2182|picorv32_core/reg25_b16  (
    .a({\picorv32_core/n669_lutinv_placeOpt_2 ,_al_u2182_o}),
    .b({\picorv32_core/mem_do_rdata ,_al_u2183_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_2 ,_al_u2184_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o_placeOpt_2,_al_u2181_o}),
    .e({\picorv32_core/pcpi_rs1$16$ ,_al_u2190_o}),
    .f({_al_u2182_o,open_n13894}),
    .q({open_n13898,\picorv32_core/pcpi_rs1$16$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(C*~(~1*~B*~(A*~D)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2184 (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .b({\picorv32_core/n576 [16],\picorv32_core/n576 [16]}),
    .c({\picorv32_core/n668_lutinv ,\picorv32_core/n668_lutinv }),
    .d({_al_u1546_o_placeOpt_2,_al_u1546_o_placeOpt_2}),
    .mi({open_n13911,\picorv32_core/mem_do_wdata }),
    .fx({open_n13916,_al_u2184_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(D*~(~A*~(1*B*~C)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010111000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2186 (
    .a({_al_u2185_o,_al_u2185_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv }),
    .c({\picorv32_core/instr_lui ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/n664_lutinv ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n13931,\picorv32_core/reg_pc [16]}),
    .fx({open_n13936,\picorv32_core/sel41_b16/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b0000001010100010),
    .MODE("LOGIC"))
    \_al_u2188|_al_u2242  (
    .a({\picorv32_core/n554 ,\picorv32_core/n554 }),
    .b({\picorv32_core/pcpi_rs1$12$ ,_al_u1302_o}),
    .c({_al_u1302_o,\picorv32_core/pcpi_rs1$10$ }),
    .d({\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/pcpi_rs1$12$ }),
    .f({_al_u2188_o,_al_u2242_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUT1("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2189 (
    .a({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .b({_al_u2187_o,_al_u2187_o}),
    .c({_al_u2188_o,_al_u2188_o}),
    .d({_al_u1313_o,_al_u1313_o}),
    .mi({open_n13971,\picorv32_core/pcpi_rs1$16$ }),
    .fx({open_n13976,\picorv32_core/sel41_b16/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*~C*~A+D*~B*~C*~A+~D*~B*~C*A+D*~B*~C*A"),
    //.LUTF1("~C*~A*~B*~D+C*~A*~B*~D+~C*~A*B*~D+C*~A*B*~D+~C*~A*B*D+C*~A*B*D"),
    //.LUTG0("D*~B*~C*~A+D*~B*~C*A"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000001100000011),
    .INIT_LUTF1(16'b0100010001010101),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2190|_al_u2234  (
    .a({\picorv32_core/sel41_b16/B5 ,open_n13979}),
    .b({_al_u1924_o,\picorv32_core/sel41_b12/B5 }),
    .c({open_n13980,\picorv32_core/sel41_b12/B2 }),
    .d({\picorv32_core/pcpi_rs1$16$ ,_al_u1924_o}),
    .e({\picorv32_core/sel41_b16/B2 ,\picorv32_core/pcpi_rs1$12$ }),
    .f({_al_u2190_o,_al_u2234_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~C*~B*~D*~A+~C*~B*~D*A"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~C*~B*~D*~A+~C*~B*D*~A+~C*~B*~D*A+~C*~B*D*A"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2192|_al_u2195  (
    .a({open_n14003,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .b({\picorv32_core/n576 [15],\picorv32_core/n576 [15]}),
    .c({\picorv32_core/mem_do_rdata ,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/mem_do_prefetch_placeOpt_2 ,_al_u1546_o_placeOpt_2}),
    .e({_al_u1546_o_placeOpt_2,\picorv32_core/mem_do_wdata }),
    .f({_al_u2192_o,_al_u2195_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTF1("~D*B*~A*~C+~D*~B*A*~C+~D*B*A*~C+~D*B*~A*C+~D*~B*A*C+~D*B*A*C"),
    //.LUTG0("(B*~(~1*~(~A*~(C*~D))))"),
    //.LUTG1("~D*~B*A*~C+~D*B*A*~C+~D*~B*A*C+~D*B*A*C"),
    .INIT_LUTF0(16'b0100010000000100),
    .INIT_LUTF1(16'b0000000011101110),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b0000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2194|_al_u2193  (
    .a({\picorv32_core/mem_do_wdata ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_2 ,\picorv32_core/n669_lutinv_placeOpt_2 }),
    .c({open_n14026,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .d({\picorv32_core/pcpi_rs1$15$ ,_al_u1546_o_placeOpt_2}),
    .e({_al_u1546_o_placeOpt_2,\picorv32_core/pcpi_rs1$15$ }),
    .f({_al_u2194_o,_al_u2193_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(C*~(~A*~(1*B*~D)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010000011100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2197 (
    .a({_al_u2196_o,_al_u2196_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv_placeOpt_2 }),
    .c({\picorv32_core/n664_lutinv_placeOpt_2 ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/instr_lui ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n14061,\picorv32_core/reg_pc [15]}),
    .fx({open_n14066,\picorv32_core/sel41_b15/B5 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+~A*B*~C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*B*C*D"),
    //.LUTF1("~B*~C*~A*~D+~B*C*~A*~D+~B*~C*A*~D+~B*C*A*~D+~B*~C*~A*D+~B*~C*A*D"),
    //.LUTG0("~A*~B*~C*~D+~A*~B*~C*D"),
    //.LUTG1("~B*C*~A*~D+~B*C*A*~D"),
    .INIT_LUTF0(16'b0100010101000101),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000000100000001),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2198|_al_u2220  (
    .a({open_n14069,\picorv32_core/n554 }),
    .b({\picorv32_core/n554 ,_al_u1302_o}),
    .c({_al_u1302_o,\picorv32_core/pcpi_rs1$12$ }),
    .d({\picorv32_core/pcpi_rs1$16$ ,open_n14072}),
    .e({\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$14$ }),
    .f({_al_u2198_o,_al_u2220_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("D*~A*~B*~C+D*A*~B*~C+D*~A*B*~C+D*A*B*~C"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("D*~A*~B*~C+D*A*~B*~C+D*~A*~B*C+D*A*~B*C"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0011001100000000),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2199|_al_u1952  (
    .b({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$11$ }),
    .c({\picorv32_core/pcpi_rs1$11$ ,\picorv32_core/pcpi_rs1$3$ }),
    .d({_al_u1302_o,\picorv32_core/n554 }),
    .e({\picorv32_core/pcpi_rs1$19$ ,_al_u1302_o}),
    .f({_al_u2199_o,_al_u1952_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    //.LUTG0("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b1010101000000010),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2201|_al_u2200  (
    .a({open_n14117,\picorv32_core/n667_lutinv }),
    .b({\picorv32_core/sel41_b15/B5 ,_al_u2198_o}),
    .c({_al_u1924_o,_al_u2199_o}),
    .d({\picorv32_core/sel41_b15/B2 ,_al_u1313_o}),
    .e({\picorv32_core/pcpi_rs1$15$ ,\picorv32_core/pcpi_rs1$15$ }),
    .f({_al_u2201_o,\picorv32_core/sel41_b15/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2203|_al_u2206  (
    .a({open_n14140,\picorv32_core/mem_do_prefetch_placeOpt_6 }),
    .b({\picorv32_core/n576 [14],\picorv32_core/n576 [14]}),
    .c({_al_u1546_o_placeOpt_8,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/mem_do_rdata ,_al_u1546_o_placeOpt_8}),
    .e({\picorv32_core/mem_do_prefetch_placeOpt_6 ,\picorv32_core/mem_do_wdata }),
    .f({_al_u2203_o,_al_u2206_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTF1("~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG0("(B*~(~1*~(~A*~(C*~D))))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0100010000000100),
    .INIT_LUTF1(16'b1111000011111010),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2205|_al_u2204  (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_6 ,\picorv32_core/mem_do_rdata }),
    .b({open_n14163,\picorv32_core/n669_lutinv_placeOpt_3 }),
    .c({\picorv32_core/mem_do_wdata ,\picorv32_core/mem_do_prefetch_placeOpt_6 }),
    .d({_al_u1546_o_placeOpt_8,_al_u1546_o_placeOpt_8}),
    .e({\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$14$ }),
    .f({_al_u2205_o,_al_u2204_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*((~C*~D)*~(0)*~(B)+(~C*~D)*0*~(B)+~((~C*~D))*0*B+(~C*~D)*0*B))"),
    //.LUTF1("~B*~C*~D*~A+B*~C*~D*~A+~B*~C*~D*A+B*~C*~D*A"),
    //.LUTG0("(A*((~C*~D)*~(1)*~(B)+(~C*~D)*1*~(B)+~((~C*~D))*1*B+(~C*~D)*1*B))"),
    //.LUTG1("~B*~C*~D*~A+B*~C*~D*~A+~B*~C*D*~A+B*~C*D*~A"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1000100010001010),
    .INIT_LUTG1(16'b0000010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2209|_al_u2211  (
    .a({\picorv32_core/pcpi_rs1$15$ ,\picorv32_core/n667_lutinv }),
    .b({open_n14186,_al_u1313_o}),
    .c({\picorv32_core/n554 ,_al_u2210_o}),
    .d({\picorv32_core/pcpi_rs1$13$ ,_al_u2209_o}),
    .e({_al_u1302_o,\picorv32_core/pcpi_rs1$14$ }),
    .f({_al_u2209_o,\picorv32_core/sel41_b14/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D"),
    //.LUTF1("0"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D+A*~B*~C*D+A*B*~C*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D"),
    .INIT_LUTF0(16'b0000000010101010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000101000001010),
    .INIT_LUTG1(16'b0000010110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2210|_al_u1963  (
    .a({_al_u1302_o,\picorv32_core/n554 }),
    .c({\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$10$ }),
    .d({\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$2$ }),
    .e({\picorv32_core/n554 ,_al_u1302_o}),
    .f({_al_u2210_o,_al_u1963_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("~B*A*~C*~D+B*A*~C*~D"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0000000000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2212|_al_u2208  (
    .a({_al_u1924_o,_al_u2207_o}),
    .b({open_n14233,\picorv32_core/n664_lutinv_placeOpt_2 }),
    .c({\picorv32_core/sel41_b14/B2 ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/sel41_b14/B5 ,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/reg_pc [14]}),
    .f({_al_u2212_o,\picorv32_core/sel41_b14/B5 }));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(D*~C)*~(B*~A))"),
    //.LUTF1("(A*~(~0*~(~B*~(C*~D))))"),
    //.LUTG0("~(1*~(D*~C)*~(B*~A))"),
    //.LUTG1("(A*~(~1*~(~B*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0010001000000010),
    .INIT_LUTG0(16'b0100111101000100),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2215|picorv32_core/reg25_b13  (
    .a({\picorv32_core/n669_lutinv_placeOpt_2 ,_al_u2214_o}),
    .b({\picorv32_core/mem_do_rdata ,_al_u2215_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_7 ,_al_u2216_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o_placeOpt_7,_al_u2217_o}),
    .e({\picorv32_core/pcpi_rs1$13$ ,_al_u2223_o}),
    .f({_al_u2215_o,open_n14271}),
    .q({open_n14275,\picorv32_core/pcpi_rs1$13$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(B*~(~1*~A*~(D*~C)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1100110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2217 (
    .a({\picorv32_core/n576 [13],\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .b({\picorv32_core/n668_lutinv ,\picorv32_core/n576 [13]}),
    .c({_al_u1546_o_placeOpt_7,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/mem_do_prefetch_placeOpt_7 ,_al_u1546_o_placeOpt_7}),
    .mi({open_n14288,\picorv32_core/mem_do_wdata }),
    .fx({open_n14293,_al_u2217_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT_LUT0(16'b0000001010001010),
    .INIT_LUT1(16'b0010000000101010),
    .MODE("LOGIC"))
    \_al_u2221|_al_u1974  (
    .a({\picorv32_core/n554 ,\picorv32_core/n554 }),
    .b({\picorv32_core/pcpi_rs1$17$ ,_al_u1302_o}),
    .c({_al_u1302_o,\picorv32_core/pcpi_rs1$1$ }),
    .d({\picorv32_core/pcpi_rs1$9$ ,\picorv32_core/pcpi_rs1$9$ }),
    .f({_al_u2221_o,_al_u1974_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUT1("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2222 (
    .a({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .b({_al_u2220_o,_al_u2220_o}),
    .c({_al_u2221_o,_al_u2221_o}),
    .d({_al_u1313_o,_al_u1313_o}),
    .mi({open_n14328,\picorv32_core/pcpi_rs1$13$ }),
    .fx({open_n14333,\picorv32_core/sel41_b13/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("~A*~B*C*~D+~A*~B*C*D"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0001000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2223|_al_u2219  (
    .a({\picorv32_core/sel41_b13/B5 ,_al_u2218_o}),
    .b({\picorv32_core/sel41_b13/B2 ,\picorv32_core/n664_lutinv_placeOpt_1 }),
    .c({_al_u1924_o,\picorv32_core/instr_lui }),
    .d({open_n14338,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/reg_pc [13]}),
    .f({_al_u2223_o,\picorv32_core/sel41_b13/B5 }));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(D*~B)*~(A*~C))"),
    //.LUTF1("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTG0("~(1*~(D*~B)*~(A*~C))"),
    //.LUTG1("(B*~(~1*~(~A*~(C*~D))))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0100010000000100),
    .INIT_LUTG0(16'b0011101100001010),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2226|picorv32_core/reg25_b12  (
    .a({\picorv32_core/mem_do_rdata ,_al_u2226_o}),
    .b({\picorv32_core/n669_lutinv_placeOpt_2 ,_al_u2227_o}),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_2 ,_al_u2225_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1546_o_placeOpt_2,_al_u2228_o}),
    .e({\picorv32_core/pcpi_rs1$12$ ,_al_u2234_o}),
    .f({_al_u2226_o,open_n14374}),
    .q({open_n14378,\picorv32_core/pcpi_rs1$12$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~B*~(A*~D)))"),
    //.LUT1("(B*~(~1*~A*~(D*~C)))"),
    .INIT_LUT0(16'b1100000011100000),
    .INIT_LUT1(16'b1100110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2228 (
    .a({\picorv32_core/n576 [12],\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .b({\picorv32_core/n668_lutinv ,\picorv32_core/n576 [12]}),
    .c({_al_u1546_o_placeOpt_7,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/mem_do_prefetch_placeOpt_2 ,_al_u1546_o_placeOpt_7}),
    .mi({open_n14391,\picorv32_core/mem_do_wdata }),
    .fx({open_n14396,_al_u2228_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(C*~(~A*~(1*B*~D)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010000011100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2230 (
    .a({_al_u2229_o,_al_u2229_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv }),
    .c({\picorv32_core/n664_lutinv ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/instr_lui ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n14411,\picorv32_core/reg_pc [12]}),
    .fx({open_n14416,\picorv32_core/sel41_b12/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT_LUT0(16'b0000010000010101),
    .INIT_LUT1(16'b0001000000010101),
    .MODE("LOGIC"))
    \_al_u2231|_al_u2253  (
    .a({\picorv32_core/n554 ,\picorv32_core/n554 }),
    .b({\picorv32_core/pcpi_rs1$13$ ,_al_u1302_o}),
    .c({_al_u1302_o,\picorv32_core/pcpi_rs1$11$ }),
    .d({\picorv32_core/pcpi_rs1$11$ ,\picorv32_core/pcpi_rs1$9$ }),
    .f({_al_u2231_o,_al_u2253_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("C*~D*~B*~A+C*D*~B*~A+C*D*B*~A+C*~D*~B*A+C*D*~B*A+C*D*B*A"),
    //.LUTF1("B*~D*~C*~A+B*D*~C*~A+B*~D*C*~A+B*~D*~C*A+B*D*~C*A+B*~D*C*A"),
    //.LUTG0("C*~D*~B*~A+C*~D*~B*A"),
    //.LUTG1("B*D*~C*~A+B*D*~C*A"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2232|_al_u1985  (
    .b({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$0$ }),
    .c({\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/n554 }),
    .d({_al_u1302_o,_al_u1302_o}),
    .e({\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/pcpi_rs1$8$ }),
    .f({_al_u2232_o,_al_u1985_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUT1("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2233 (
    .a({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .b({_al_u2231_o,_al_u2231_o}),
    .c({_al_u2232_o,_al_u2232_o}),
    .d({_al_u1313_o,_al_u1313_o}),
    .mi({open_n14475,\picorv32_core/pcpi_rs1$12$ }),
    .fx({open_n14480,\picorv32_core/sel41_b12/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~C*~D*~B*~A+~C*~D*~B*A"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~C*~D*~B*~A+~C*~D*B*~A+~C*~D*~B*A+~C*~D*B*A"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2236|_al_u2239  (
    .a({open_n14483,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_7 ,\picorv32_core/n576 [11]}),
    .c({\picorv32_core/mem_do_rdata ,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/n576 [11],_al_u1546_o_placeOpt_7}),
    .e({_al_u1546_o_placeOpt_7,\picorv32_core/mem_do_wdata }),
    .f({_al_u2236_o,_al_u2239_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUT1("(C*~(~1*~(~B*~(A*~D))))"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b1111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2237 (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_7 ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_rdata ,\picorv32_core/n669_lutinv_placeOpt_2 }),
    .c({\picorv32_core/n669_lutinv_placeOpt_2 ,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .d({_al_u1546_o_placeOpt_7,_al_u1546_o_placeOpt_7}),
    .mi({open_n14518,\picorv32_core/pcpi_rs1$11$ }),
    .fx({open_n14523,_al_u2237_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(D*~(~A*~(1*B*~C)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010111000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2241 (
    .a({_al_u2240_o,_al_u2240_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv_placeOpt_2 }),
    .c({\picorv32_core/instr_lui ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/n664_lutinv_placeOpt_2 ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n14538,\picorv32_core/reg_pc [11]}),
    .fx({open_n14543,\picorv32_core/sel41_b11/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*~(B*~D)))"),
    //.LUT1("(A*~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUT0(16'b0101000001010100),
    .INIT_LUT1(16'b0000101000100010),
    .MODE("LOGIC"))
    \_al_u2243|_al_u1947  (
    .a({\picorv32_core/n554 ,\picorv32_core/pcpi_rs1$7$ }),
    .b({\picorv32_core/pcpi_rs1$7$ ,\picorv32_core/mem_do_prefetch_placeOpt_2 }),
    .c({\picorv32_core/pcpi_rs1$15$ ,\picorv32_core/mem_do_wdata }),
    .d({_al_u1302_o,_al_u1546_o_placeOpt_2}),
    .f({_al_u2243_o,_al_u1947_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUTF1("~B*~A*~C*~D+~B*A*~C*~D+~B*~A*C*~D+~B*A*C*~D"),
    //.LUTG0("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    //.LUTG1("~B*~A*C*~D+~B*A*C*~D"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b1010101000000010),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2245|_al_u2244  (
    .a({open_n14566,\picorv32_core/n667_lutinv }),
    .b({\picorv32_core/sel41_b11/B5 ,_al_u2242_o}),
    .c({_al_u1924_o,_al_u2243_o}),
    .d({\picorv32_core/sel41_b11/B2 ,_al_u1313_o}),
    .e({\picorv32_core/pcpi_rs1$11$ ,\picorv32_core/pcpi_rs1$11$ }),
    .f({_al_u2245_o,\picorv32_core/sel41_b11/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~0*~B*~(A*~D)))"),
    //.LUTF1("~A*~B*~C*~D+~A*~B*C*~D"),
    //.LUTG0("(C*~(~1*~B*~(A*~D)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000000000010001),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2247|_al_u2250  (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_4 ,\picorv32_core/mem_do_prefetch_placeOpt_4 }),
    .b({\picorv32_core/n576 [10],\picorv32_core/n576 [10]}),
    .c({open_n14589,\picorv32_core/n668_lutinv }),
    .d({\picorv32_core/mem_do_rdata ,_al_u1546_o_placeOpt_5}),
    .e({_al_u1546_o_placeOpt_5,\picorv32_core/mem_do_wdata }),
    .f({_al_u2247_o,_al_u2250_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUTF1("~A*B*~D*~C+~A*~B*D*~C+~A*B*D*~C+~A*B*~D*C+~A*~B*D*C+~A*B*D*C"),
    //.LUTG0("(B*~(~1*~(~A*~(C*~D))))"),
    //.LUTG1("~A*~B*D*~C+~A*B*D*~C+~A*~B*D*C+~A*B*D*C"),
    .INIT_LUTF0(16'b0100010000000100),
    .INIT_LUTF1(16'b0101010101000100),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b0101010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2249|_al_u2248  (
    .a({\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/mem_do_prefetch_placeOpt_4 ,\picorv32_core/n669_lutinv_placeOpt_3 }),
    .c({open_n14612,\picorv32_core/mem_do_prefetch_placeOpt_4 }),
    .d({\picorv32_core/mem_do_wdata ,_al_u1546_o_placeOpt_5}),
    .e({_al_u1546_o_placeOpt_5,\picorv32_core/pcpi_rs1$10$ }),
    .f({_al_u2249_o,_al_u2248_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*((~C*~B)*~(0)*~(D)+(~C*~B)*0*~(D)+~((~C*~B))*0*D+(~C*~B)*0*D))"),
    //.LUT1("(A*((~C*~B)*~(1)*~(D)+(~C*~B)*1*~(D)+~((~C*~B))*1*D+(~C*~B)*1*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2255 (
    .a({\picorv32_core/n667_lutinv ,\picorv32_core/n667_lutinv }),
    .b({_al_u2253_o,_al_u2253_o}),
    .c({_al_u2254_o,_al_u2254_o}),
    .d({_al_u1313_o,_al_u1313_o}),
    .mi({open_n14647,\picorv32_core/pcpi_rs1$10$ }),
    .fx({open_n14652,\picorv32_core/sel41_b10/B2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(0*D*~C)))"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D"),
    //.LUTG0("(B*~(~A*~(1*D*~C)))"),
    //.LUTG1("~B*A*~C*~D+B*A*~C*~D"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b0000000000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2256|_al_u2252  (
    .a({_al_u1924_o,_al_u2251_o}),
    .b({open_n14655,\picorv32_core/n664_lutinv_placeOpt_4 }),
    .c({\picorv32_core/sel41_b10/B2 ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/sel41_b10/B5 ,\picorv32_core/is_lui_auipc_jal }),
    .e({\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/reg_pc [10]}),
    .f({_al_u2256_o,\picorv32_core/sel41_b10/B5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~0*~(~A*~(C*~D))))"),
    //.LUT1("(B*~(~1*~(~A*~(C*~D))))"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b1100110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2259 (
    .a({\picorv32_core/mem_do_rdata ,\picorv32_core/mem_do_rdata }),
    .b({\picorv32_core/n669_lutinv_placeOpt_4 ,\picorv32_core/n669_lutinv_placeOpt_4 }),
    .c({\picorv32_core/mem_do_prefetch_placeOpt_8 ,\picorv32_core/mem_do_prefetch_placeOpt_8 }),
    .d({_al_u1546_o_placeOpt_8,_al_u1546_o_placeOpt_8}),
    .mi({open_n14690,\picorv32_core/pcpi_rs1$0$ }),
    .fx({open_n14695,_al_u2259_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~0*~C*~(A*~D)))"),
    //.LUT1("(B*~(~1*~C*~(A*~D)))"),
    .INIT_LUT0(16'b1100000011001000),
    .INIT_LUT1(16'b1100110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2261 (
    .a({\picorv32_core/mem_do_prefetch_placeOpt_8 ,\picorv32_core/mem_do_prefetch_placeOpt_8 }),
    .b({\picorv32_core/n668_lutinv ,\picorv32_core/n668_lutinv }),
    .c({\picorv32_core/n576 [0],\picorv32_core/n576 [0]}),
    .d({_al_u1546_o_placeOpt_8,_al_u1546_o_placeOpt_8}),
    .mi({open_n14710,\picorv32_core/mem_do_wdata }),
    .fx({open_n14715,_al_u2261_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*A*(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B))"),
    //.LUT1("(C*A*(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B))"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b1010000010000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2262 (
    .a({\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv ,\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv }),
    .b({\picorv32_core/n554 ,\picorv32_core/n554 }),
    .c({_al_u1302_o,_al_u1302_o}),
    .d({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$1$ }),
    .mi({open_n14730,\picorv32_core/pcpi_rs1$4$ }),
    .fx({open_n14735,_al_u2262_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(0*D*~C)))"),
    //.LUT1("(D*~(~A*~(1*B*~C)))"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010111000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2264 (
    .a({_al_u2263_o,_al_u2263_o}),
    .b({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/n664_lutinv_placeOpt_3 }),
    .c({\picorv32_core/instr_lui ,\picorv32_core/instr_lui }),
    .d({\picorv32_core/n664_lutinv_placeOpt_3 ,\picorv32_core/is_lui_auipc_jal }),
    .mi({open_n14750,\picorv32_core/reg_pc [0]}),
    .fx({open_n14755,\picorv32_core/sel41_b0/B5 }));
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~((A*D))+B*C*~((A*D))+~(B)*C*(A*D)+B*C*(A*D))"),
    //.LUT1("~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110010011001100),
    .INIT_LUT1(16'b0000101001011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2268|picorv32_core/reg6_b1  (
    .a({\picorv32_core/mem_xfer ,\picorv32_core/mem_rdata_latched [0]}),
    .b({open_n14758,\picorv32_core/mem_rdata_latched [3]}),
    .c({\picorv32_core/mem_rdata_latched [21],\picorv32_core/mem_rdata_latched [21]}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [21],\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .f({_al_u2268_o,open_n14772}),
    .q({open_n14776,\picorv32_core/decoded_imm_uj [1]}));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~A*~(D*~(~0*~C)))"),
    //.LUTF1("(~B*C*~(D*~(~0*~A)))"),
    //.LUTG0("(~B*~A*~(D*~(~1*~C)))"),
    //.LUTG1("(~B*C*~(D*~(~1*~A)))"),
    .INIT_LUTF0(16'b0000000100010001),
    .INIT_LUTF1(16'b0001000000110000),
    .INIT_LUTG0(16'b0000000000010001),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2271|_al_u1625  (
    .a({_al_u1431_o,_al_u1481_o}),
    .b({_al_u1538_o,_al_u1538_o}),
    .c({\picorv32_core/mem_rdata_latched [12],_al_u1431_o}),
    .d({_al_u1537_o,_al_u1537_o}),
    .e({_al_u1088_o,_al_u1088_o}),
    .f({_al_u2271_o,_al_u1625_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(0*C*~(B*D*A))"),
    //.LUT1("(1*C*~(B*D*A))"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2272 (
    .a({_al_u1634_o,_al_u1634_o}),
    .b({\picorv32_core/mux79_b1/B0_3 ,\picorv32_core/mux79_b1/B0_3 }),
    .c({_al_u2271_o,_al_u2271_o}),
    .d({_al_u2270_o,_al_u2270_o}),
    .mi({open_n14811,_al_u1485_o_placeOpt_1}),
    .fx({open_n14816,_al_u2272_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*D*C*A+B*D*C*A"),
    //.LUTF1("C*~A*~D*B+C*A*~D*B"),
    //.LUTG0("~B*~D*C*A+B*~D*C*A+~B*D*C*A+B*D*C*A"),
    //.LUTG1("~C*~A*~D*B+C*~A*~D*B+~C*A*~D*B+C*A*~D*B"),
    .INIT_LUTF0(16'b1010000000000000),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b1010000010100000),
    .INIT_LUTG1(16'b0000000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2273|_al_u2460  (
    .a({open_n14819,_al_u1546_o}),
    .b({_al_u1546_o,open_n14820}),
    .c({\picorv32_core/mem_do_prefetch ,\picorv32_core/mem_rdata_latched$0$_placeOpt_2 }),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_3 ,\picorv32_core/mem_do_prefetch }),
    .e({\picorv32_core/mem_do_rinst ,\picorv32_core/mem_do_rinst }),
    .f({_al_u2273_o,_al_u2460_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(A*~((~B*~D))*~(0)+A*(~B*~D)*~(0)+~(A)*(~B*~D)*0+A*(~B*~D)*0))"),
    //.LUT1("(~A*~(D*~((~B*~C))*~(1)+D*(~B*~C)*~(1)+~(D)*(~B*~C)*1+D*(~B*~C)*1))"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b0101010001010100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2275 (
    .a({_al_u1481_o_placeOpt_2,\picorv32_core/mem_rdata_latched [3]}),
    .b({_al_u1483_o_placeOpt_2,_al_u1483_o_placeOpt_2}),
    .c({_al_u2268_o,_al_u1481_o_placeOpt_2}),
    .d({\picorv32_core/mem_rdata_latched [3],_al_u2268_o}),
    .mi({open_n14855,_al_u1485_o_placeOpt_3}),
    .fx({open_n14860,_al_u2275_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D)))"),
    //.LUTF1("(C*~(~B*~(A*~(0*~D))))"),
    //.LUTG0("(A*~(1*~(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D)))"),
    //.LUTG1("(C*~(~B*~(A*~(1*~D))))"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b1110000011100000),
    .INIT_LUTG0(16'b1000100000001010),
    .INIT_LUTG1(16'b1110000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2276|_al_u2269  (
    .a({_al_u2269_o,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .b({_al_u2274_o,\picorv32_core/mem_rdata_latched [3]}),
    .c({_al_u2273_o,_al_u2268_o}),
    .d({_al_u2272_o,_al_u2267_o}),
    .e({_al_u2275_o,_al_u1481_o_placeOpt_2}),
    .f({_al_u2276_o,_al_u2269_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~A*~B*C*D)"),
    //.LUT1("(~1*~A*~B*C*D)"),
    .INIT_LUT0(16'b0001000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2277 (
    .a({\picorv32_core/mem_rdata_latched [3],\picorv32_core/mem_rdata_latched [3]}),
    .b({\picorv32_core/mem_rdata_latched [4],\picorv32_core/mem_rdata_latched [4]}),
    .c({_al_u1498_o,_al_u1498_o}),
    .d({\picorv32_core/n98_lutinv ,\picorv32_core/n98_lutinv }),
    .mi({open_n14897,\picorv32_core/mem_rdata_latched [2]}),
    .fx({open_n14902,_al_u2277_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~0*~(~B*~(~C*D))))"),
    //.LUT1("(B*~(~1*~(~A*~(~C*D))))"),
    .INIT_LUT0(16'b0010000000100010),
    .INIT_LUT1(16'b1100110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2279 (
    .a({_al_u2278_o,\picorv32_core/mem_rdata_latched$1$_placeOpt_1 }),
    .b({\picorv32_core/mem_rdata_latched$1$_placeOpt_1 ,_al_u2278_o}),
    .c({_al_u1635_o,_al_u1635_o}),
    .d({_al_u2277_o,_al_u2277_o}),
    .mi({open_n14917,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .fx({open_n14922,_al_u2279_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D"),
    //.LUTG1("A*~B*~C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b0000000000001010),
    .INIT_LUTF1(16'b0111011101110111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0010001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2281|_al_u2283  (
    .a({\picorv32_core/mem_xfer ,_al_u1485_o_placeOpt_3}),
    .b({\picorv32_core/mem_rdata_latched [20],open_n14925}),
    .c({open_n14926,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .d({open_n14929,_al_u2281_o}),
    .e({\picorv32_core/mem_rdata_q [20],_al_u1481_o_placeOpt_4}),
    .f({_al_u2281_o,_al_u2283_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(A*~((~C*~D))*~(0)+A*(~C*~D)*~(0)+~(A)*(~C*~D)*0+A*(~C*~D)*0))"),
    //.LUT1("(~A*~(D*~((~B*~C))*~(1)+D*(~B*~C)*~(1)+~(D)*(~B*~C)*1+D*(~B*~C)*1))"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0101010001010100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2284 (
    .a({_al_u1481_o_placeOpt_2,\picorv32_core/mem_rdata_latched [2]}),
    .b({_al_u1483_o_placeOpt_2,_al_u1481_o_placeOpt_2}),
    .c({_al_u2281_o,_al_u1483_o_placeOpt_2}),
    .d({\picorv32_core/mem_rdata_latched [2],_al_u2281_o}),
    .mi({open_n14962,_al_u1485_o_placeOpt_3}),
    .fx({open_n14967,_al_u2284_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)))"),
    //.LUTF1("(C*~(~B*~(A*~(0*~D))))"),
    //.LUTG0("(A*~(1*~(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)))"),
    //.LUTG1("(C*~(~B*~(A*~(1*~D))))"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b1110000011100000),
    .INIT_LUTG0(16'b1000000010100010),
    .INIT_LUTG1(16'b1110000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2285|_al_u2282  (
    .a({_al_u2282_o,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .b({_al_u2283_o,_al_u2267_o}),
    .c({_al_u2273_o,\picorv32_core/mem_rdata_latched [2]}),
    .d({_al_u2272_o,_al_u2281_o}),
    .e({_al_u2284_o,_al_u1481_o_placeOpt_2}),
    .f({_al_u2285_o,_al_u2282_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(0*~A*~B*~C*D)"),
    //.LUT1("(1*~B*~A*~C*D)"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2287 (
    .a(\picorv32_core/mem_rdata_latched [3:2]),
    .b({\picorv32_core/mem_rdata_latched [2],\picorv32_core/mem_rdata_latched [3]}),
    .c({\picorv32_core/mem_rdata_latched [4],\picorv32_core/mem_rdata_latched [4]}),
    .d({_al_u1498_o,_al_u1498_o}),
    .mi({open_n15004,\picorv32_core/mem_rdata_latched [12]}),
    .fx({open_n15009,_al_u2287_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(~A*~B*~C*D))"),
    //.LUT1("(1*~(~B*~A*~C*D))"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1111111011111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2288 (
    .a(\picorv32_core/mem_rdata_latched [3:2]),
    .b({\picorv32_core/mem_rdata_latched [2],\picorv32_core/mem_rdata_latched [3]}),
    .c({\picorv32_core/mem_rdata_latched [4],\picorv32_core/mem_rdata_latched [4]}),
    .d({_al_u1498_o,_al_u1498_o}),
    .mi({open_n15024,\picorv32_core/mux79_b0/B0_3 }),
    .fx({open_n15029,_al_u2288_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*~A)"),
    //.LUTF1("(~0*~(A*~(~C*~(~B*D))))"),
    //.LUTG0("(~1*~D*~C*~B*~A)"),
    //.LUTG1("(~1*~(A*~(~C*~(~B*D))))"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0101110101011111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2290|_al_u1654  (
    .a({\picorv32_core/n98_lutinv ,\picorv32_core/mux79_b1/B0_3 }),
    .b({_al_u1654_o,_al_u1444_o}),
    .c({_al_u2288_o,\picorv32_core/mux79_b2/B0_3 }),
    .d({_al_u2287_o,\picorv32_core/mux79_b0/B0_3 }),
    .e({_al_u2289_o,_al_u1464_o}),
    .f({_al_u2290_o,_al_u1654_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*C*D)"),
    //.LUT1("(B*A*D)"),
    .INIT_LUT0(16'b0101000000000000),
    .INIT_LUT1(16'b1000100000000000),
    .MODE("LOGIC"))
    \_al_u2295|_al_u1630  (
    .a({_al_u1444_o,_al_u1464_o}),
    .b({_al_u1464_o,open_n15054}),
    .c({open_n15055,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .d({\picorv32_core/mem_rdata_latched [12],\picorv32_core/mem_rdata_latched [6]}),
    .f({_al_u2295_o,_al_u1630_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000001010101),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2296|_al_u2289  (
    .a({_al_u1485_o_placeOpt_3,_al_u1485_o_placeOpt_3}),
    .d({open_n15082,_al_u1481_o_placeOpt_2}),
    .e({\picorv32_core/mux79_b0/B0_3 ,\picorv32_core/mux79_b0/B0_3 }),
    .f({_al_u2296_o,_al_u2289_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~B)"),
    //.LUT1("(~B*C*A*~D)"),
    .INIT_LUT0(16'b0011001100000000),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"))
    \_al_u2297|_al_u1536  (
    .a({_al_u1536_o,open_n15103}),
    .b({_al_u1483_o_placeOpt_2,\picorv32_core/mem_rdata_latched$1$_placeOpt_1 }),
    .c({_al_u2296_o,open_n15104}),
    .d({_al_u2295_o,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .f({_al_u2297_o,_al_u1536_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~C*~(~A*D))"),
    //.LUT1("(B*~(D*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011111110011),
    .INIT_LUT1(16'b1000100011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2300|picorv32_core/reg22_b6  (
    .a({_al_u1546_o_placeOpt_1,_al_u1184_o}),
    .b({\picorv32_core/n666_lutinv ,_al_u2302_o}),
    .c({open_n15125,\picorv32_core/sel40_b6/B3 }),
    .clk(clk_pad),
    .d({\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ,\picorv32_core/n580 }),
    .sr(\picorv32_core/mux164_b0_sel_is_0_o ),
    .f({\picorv32_core/sel40_b6/B3 ,open_n15139}),
    .q({open_n15143,\picorv32_core/cpu_state [6]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~A*~(C*B))"),
    //.LUT1("(~B*A)"),
    .INIT_LUT0(16'b0001010100000000),
    .INIT_LUT1(16'b0010001000100010),
    .MODE("LOGIC"))
    \_al_u2302|_al_u2301  (
    .a({_al_u2301_o,\picorv32_core/sel40_b6/B5 }),
    .b({_al_u1550_o,\picorv32_core/n667_lutinv }),
    .c({open_n15144,_al_u1313_o}),
    .d({open_n15147,resetn_placeOpt_16}),
    .f({_al_u2302_o,_al_u2301_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~0*~D*C)*~(B*~A))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTG0("(~(~1*~D*C)*~(B*~A))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1011101100001011),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b1011101110111011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2305|_al_u2306  (
    .a({\picorv32_core/n523_lutinv ,_al_u2305_o}),
    .b({\picorv32_core/is_sll_srl_sra ,\picorv32_core/n664_lutinv_placeOpt_2 }),
    .c({\picorv32_core/is_jalr_addi_slti_sltiu_xori_ori_andi ,\picorv32_core/n665_lutinv }),
    .d({\picorv32_core/is_sb_sh_sw ,\picorv32_core/is_sb_sh_sw }),
    .e({\picorv32_core/is_lui_auipc_jal ,\picorv32_core/is_sll_srl_sra }),
    .f({_al_u2305_o,_al_u2306_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0100110001001100),
    .INIT_LUTG0(16'b0101010101010101),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2307|picorv32_core/reg22_b3  (
    .a({\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ,_al_u2307_o}),
    .b({_al_u2306_o,open_n15188}),
    .c({\picorv32_core/n666_lutinv ,open_n15189}),
    .clk(clk_pad),
    .e({_al_u1546_o_placeOpt_1,resetn_placeOpt_8}),
    .sr(\picorv32_core/mux164_b0_sel_is_0_o ),
    .f({_al_u2307_o,open_n15207}),
    .q({open_n15211,\picorv32_core/cpu_state [3]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C)*~(0*B))"),
    //.LUT1("(~A*~(D*C)*~(1*B))"),
    .INIT_LUT0(16'b0000010101010101),
    .INIT_LUT1(16'b0000000100010001),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2309 (
    .a({\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv ,\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv }),
    .b({\picorv32_core/n664_lutinv_placeOpt_1 ,\picorv32_core/n664_lutinv_placeOpt_1 }),
    .c({\picorv32_core/n665_lutinv ,\picorv32_core/n665_lutinv }),
    .d({\picorv32_core/is_sll_srl_sra ,\picorv32_core/is_sll_srl_sra }),
    .mi({open_n15224,\picorv32_core/is_slli_srli_srai }),
    .fx({open_n15229,_al_u2309_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~A*C*~B*~D+~A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0101111101010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2310|picorv32_core/reg22_b2  (
    .a({\picorv32_core/is_sll_srl_sra ,open_n15232}),
    .c({\picorv32_core/n664_lutinv_placeOpt_1 ,resetn_placeOpt_8}),
    .clk(clk_pad),
    .d({_al_u2309_o,_al_u2310_o}),
    .e({\picorv32_core/n523_lutinv ,open_n15236}),
    .sr(\picorv32_core/mux164_b0_sel_is_0_o ),
    .f({_al_u2310_o,open_n15251}),
    .q({open_n15255,\picorv32_core/cpu_state [2]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(~C*~(A*~(~B*D))))"),
    //.LUTF1("~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG0("(1*~(~C*~(A*~(~B*D))))"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b1111100011111010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2312|picorv32_core/reg22_b1  (
    .a({open_n15256,\picorv32_core/n668_lutinv }),
    .b({open_n15257,\picorv32_core/mem_do_prefetch_placeOpt_7 }),
    .c({open_n15258,\picorv32_core/sel40_b1/or_or_B4_B5_o_or_B6__o_lutinv }),
    .clk(clk_pad),
    .d({\picorv32_core/is_sb_sh_sw ,_al_u1546_o_placeOpt_1}),
    .e({_al_u1337_o,resetn_placeOpt_16}),
    .sr(\picorv32_core/mux164_b0_sel_is_0_o ),
    .f({\picorv32_core/sel40_b1/or_or_B4_B5_o_or_B6__o_lutinv ,open_n15274}),
    .q({open_n15278,\picorv32_core/cpu_state [1]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*A*~B*~C+D*A*~B*~C+~D*A*B*~C+D*A*B*~C+~D*A*~B*C+D*A*~B*C+~D*A*B*C+D*A*B*C"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~D*A*~B*~C+D*A*~B*~C+~D*A*B*~C+D*A*B*~C+~D*~A*B*C+D*~A*B*C+~D*A*B*C+D*A*B*C"),
    //.LUTG1("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b1101110111011101),
    .INIT_LUTG0(16'b1100101011001010),
    .INIT_LUTG1(16'b0001000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2316|picorv32_core/reg6_b4  (
    .a({\picorv32_core/mem_rdata_q [24],_al_u1464_o}),
    .b({\picorv32_core/mem_xfer ,\picorv32_core/mem_rdata_latched [24]}),
    .c({open_n15279,\picorv32_core/mem_rdata_latched [1]}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .e({\picorv32_core/mem_rdata_latched [24],\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }),
    .f({_al_u2316_o,open_n15297}),
    .q({open_n15301,\picorv32_core/decoded_imm_uj [4]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(~C*~(D*~(0*~A))))"),
    //.LUTF1("(A*~B*~(~0*~(~D*~C)))"),
    //.LUTG0("~(~B*~(~C*~(D*~(1*~A))))"),
    //.LUTG1("(A*~B*~(~1*~(~D*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011001111),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1100110111001111),
    .INIT_LUTG1(16'b0010001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2317|picorv32_core/reg0_b24  (
    .a({\picorv32_core/mem_rdata_latched$1$_placeOpt_1 ,_al_u2324_o}),
    .b({_al_u2316_o,_al_u2317_o}),
    .c({_al_u2315_o,_al_u2325_o}),
    .clk(clk_pad),
    .d({_al_u2278_o,_al_u2321_o}),
    .e({\picorv32_core/mem_rdata_latched$0$_placeOpt_4 ,_al_u2293_o}),
    .f({_al_u2317_o,open_n15318}),
    .q({open_n15322,\picorv32_core/mem_rdata_q [24]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("(0*B*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUT1("(1*B*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1000100000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2318 (
    .a({\picorv32_core/mem_rdata_latched [6],\picorv32_core/mem_rdata_latched [6]}),
    .b({_al_u1536_o,_al_u1536_o}),
    .c({_al_u2316_o,_al_u2316_o}),
    .d({_al_u2267_o,_al_u2267_o}),
    .mi({open_n15335,_al_u1481_o_placeOpt_2}),
    .fx({open_n15340,_al_u2318_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*C*~B)"),
    //.LUTF1("0"),
    //.LUTG0("(~A*C*~B)"),
    //.LUTG1("C*~A*~B*D+C*A*~B*D"),
    .INIT_LUTF0(16'b0001000000010000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0001000000010000),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2319|_al_u2278  (
    .a({open_n15343,_al_u1485_o_placeOpt_3}),
    .b({\picorv32_core/mem_rdata_latched$0$_placeOpt_4 ,_al_u1481_o_placeOpt_2}),
    .c({\picorv32_core/mem_rdata_latched$1$_placeOpt_1 ,_al_u1483_o_placeOpt_2}),
    .d({_al_u2278_o,open_n15346}),
    .e({\picorv32_core/mem_rdata_latched [6],open_n15347}),
    .f({_al_u2319_o,_al_u2278_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(~B*~(C)*~((~0*~A))+~B*C*~((~0*~A))+~(~B)*C*(~0*~A)+~B*C*(~0*~A)))"),
    //.LUT1("(D*(~B*~(C)*~((~1*~A))+~B*C*~((~1*~A))+~(~B)*C*(~1*~A)+~B*C*(~1*~A)))"),
    .INIT_LUT0(16'b0111001000000000),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2320 (
    .a({_al_u1481_o_placeOpt_2,_al_u1481_o_placeOpt_2}),
    .b({_al_u2316_o,_al_u2316_o}),
    .c({_al_u1464_o,_al_u1464_o}),
    .d({_al_u1650_o,_al_u1650_o}),
    .mi({open_n15380,_al_u1485_o_placeOpt_3}),
    .fx({open_n15385,_al_u2320_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000100000000),
    .INIT_LUTG0(16'b0011001100110011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2321|_al_u2439  (
    .a({_al_u2318_o,open_n15388}),
    .b({_al_u2319_o,_al_u1483_o_placeOpt_2}),
    .d({_al_u1569_o,open_n15393}),
    .e({_al_u2320_o,_al_u2296_o}),
    .f({_al_u2321_o,\picorv32_core/mux79_b0/B1_0 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*A*D*~(B*~C))"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D"),
    //.LUTG0("(~1*A*D*~(B*~C))"),
    //.LUTG1("B*~A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+B*~A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    .INIT_LUTF0(16'b1010001000000000),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2322|_al_u1629  (
    .a({open_n15414,\picorv32_core/mem_rdata_latched [6]}),
    .b({_al_u2316_o,_al_u1483_o_placeOpt_2}),
    .c({_al_u1483_o_placeOpt_2,_al_u1481_o_placeOpt_4}),
    .d({\picorv32_core/mem_rdata_latched [6],_al_u1606_o}),
    .e({_al_u1485_o_placeOpt_3,_al_u1485_o_placeOpt_3}),
    .f({_al_u2322_o,_al_u1629_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*~B*A*D+C*~B*A*D"),
    //.LUTF1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTG0("~C*~B*~A*~D+~C*~B*A*~D+~C*~B*~A*D+~C*~B*A*D"),
    //.LUTG1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    .INIT_LUTF0(16'b0011001100110011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000001100000011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2325|_al_u2335  (
    .b({open_n15439,_al_u2327_o}),
    .c({_al_u1569_o,_al_u1569_o}),
    .d({_al_u2316_o,open_n15442}),
    .e({open_n15443,\picorv32_core/n180 }),
    .f({_al_u2325_o,_al_u2335_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~((A*C))*~((~0*~B))+~D*(A*C)*~((~0*~B))+~(~D)*(A*C)*(~0*~B)+~D*(A*C)*(~0*~B))"),
    //.LUTF1("0"),
    //.LUTG0("~(~D*~((A*C))*~((~1*~B))+~D*(A*C)*~((~1*~B))+~(~D)*(A*C)*(~1*~B)+~D*(A*C)*(~1*~B))"),
    //.LUTG1("~B*~C*~D*~A+B*~C*~D*~A+~B*C*~D*~A+B*C*~D*~A+~B*~C*D*~A+B*~C*D*~A+~B*C*D*~A+B*C*D*~A+B*C*~D*A+B*C*D*A"),
    .INIT_LUTF0(16'b1101111100010011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1101010111010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2330|_al_u2328  (
    .a({_al_u2328_o,_al_u1483_o_placeOpt_1}),
    .b({_al_u2329_o,_al_u1481_o_placeOpt_3}),
    .c({\picorv32_core/mem_rdata_latched [5],_al_u1444_o}),
    .d({open_n15466,_al_u2327_o}),
    .e({_al_u1650_o,_al_u1485_o_placeOpt_2}),
    .f({_al_u2330_o,_al_u2328_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)))"),
    //.LUT1("(B*~(1*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D)))"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b1100000001000100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2331 (
    .a({_al_u2327_o,\picorv32_core/mem_rdata_latched [5]}),
    .b({_al_u1536_o,_al_u1536_o}),
    .c({\picorv32_core/mem_rdata_latched [5],_al_u2327_o}),
    .d({_al_u2267_o,_al_u2267_o}),
    .mi({open_n15499,_al_u1481_o_placeOpt_2}),
    .fx({open_n15504,_al_u2331_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~D*~A))"),
    //.LUTF1("~B*~D*~A*~C+~B*D*~A*~C+~B*D*A*~C+~B*~D*~A*C+~B*D*~A*C+~B*D*A*C"),
    //.LUTG0("(B*~(~D*~A))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1100110010001000),
    .INIT_LUTF1(16'b0011001100010001),
    .INIT_LUTG0(16'b1100110010001000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2332|_al_u2360  (
    .a({\picorv32_core/mux81_sel_is_1_o ,\picorv32_core/mux81_sel_is_1_o }),
    .b({_al_u1481_o_placeOpt_3,\picorv32_core/mem_rdata_latched$0$_placeOpt_1 }),
    .d({_al_u2327_o,\picorv32_core/mem_rdata_latched$1$_placeOpt_1 }),
    .e({\picorv32_core/sel10_b3/B1_1 ,open_n15511}),
    .f({_al_u2332_o,_al_u2360_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~D*~(0*A*C))"),
    //.LUTF1("~A*~C*~D*~B+~A*~C*D*~B+~A*C*D*~B+~A*~C*~D*B+~A*~C*D*B+~A*C*D*B"),
    //.LUTG0("(B*~D*~(1*A*C))"),
    //.LUTG1("~A*~C*~D*~B+~A*~C*D*~B+~A*~C*~D*B+~A*~C*D*B"),
    .INIT_LUTF0(16'b0000000011001100),
    .INIT_LUTF1(16'b0101010100000101),
    .INIT_LUTG0(16'b0000000001001100),
    .INIT_LUTG1(16'b0000010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2333|_al_u2324  (
    .a({_al_u2330_o,_al_u2323_o}),
    .b({open_n15532,_al_u2322_o}),
    .c({_al_u2331_o,_al_u1579_o}),
    .d({_al_u2332_o,_al_u2272_o}),
    .e({_al_u2272_o,\picorv32_core/mem_rdata_latched [6]}),
    .f({_al_u2333_o,_al_u2324_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D)*~(C)*~(B)*~(A)*~(0)+~(D)*C*~(B)*~(A)*~(0)+D*C*~(B)*~(A)*~(0)+~(D)*~(C)*~(B)*~(A)*0+~(D)*C*~(B)*~(A)*0+D*C*~(B)*~(A)*0+~(D)*~(C)*B*~(A)*0+~(D)*C*B*~(A)*0+D*C*B*~(A)*0+~(D)*~(C)*B*A*0+~(D)*C*B*A*0)"),
    //.LUT1("(~(D)*~(C)*~(B)*~(A)*~(1)+~(D)*C*~(B)*~(A)*~(1)+D*C*~(B)*~(A)*~(1)+~(D)*~(C)*~(B)*~(A)*1+~(D)*C*~(B)*~(A)*1+D*C*~(B)*~(A)*1+~(D)*~(C)*B*~(A)*1+~(D)*C*B*~(A)*1+D*C*B*~(A)*1+~(D)*~(C)*B*A*1+~(D)*C*B*A*1)"),
    .INIT_LUT0(16'b0001000000010001),
    .INIT_LUT1(16'b0101000011011101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2334 (
    .a({_al_u2327_o,_al_u2327_o}),
    .b({_al_u2278_o,_al_u2278_o}),
    .c({_al_u1635_o,_al_u1635_o}),
    .d({_al_u2277_o,_al_u2277_o}),
    .mi({open_n15567,\picorv32_core/mem_rdata_latched [5]}),
    .fx({open_n15572,_al_u2334_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("A*D*C*~B+A*D*C*B"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D"),
    //.LUTG0("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+~A*D*C*~B+A*D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+~A*D*C*B+A*D*C*B"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010000000000000),
    .INIT_LUTF1(16'b0000010111110101),
    .INIT_LUTG0(16'b1111111101011111),
    .INIT_LUTG1(16'b0000010111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2337|picorv32_core/reg6_b2  (
    .a({\picorv32_core/mem_rdata_q [22],\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }),
    .c({\picorv32_core/mem_xfer ,\picorv32_core/mem_rdata_latched [1]}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched [22],\picorv32_core/mem_rdata_latched [22]}),
    .e({open_n15577,\picorv32_core/mem_rdata_latched [4]}),
    .f({_al_u2337_o,open_n15593}),
    .q({open_n15597,\picorv32_core/decoded_imm_uj [2]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B*C*~A)"),
    //.LUT1("(C*~(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    .INIT_LUT0(16'b0000000000010000),
    .INIT_LUT1(16'b0111000000100000),
    .MODE("LOGIC"))
    \_al_u2338|_al_u2267  (
    .a({_al_u2267_o,_al_u1444_o}),
    .b({\picorv32_core/mem_rdata_latched [4],_al_u1483_o_placeOpt_2}),
    .c({_al_u1481_o_placeOpt_2,_al_u1464_o}),
    .d({_al_u2337_o,_al_u1485_o_placeOpt_3}),
    .f({_al_u2338_o,_al_u2267_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(A*~((~B*~D))*~(0)+A*(~B*~D)*~(0)+~(A)*(~B*~D)*0+A*(~B*~D)*0))"),
    //.LUTF1("~C*~D*~A*B+C*~D*~A*B+~C*D*~A*B+C*D*~A*B+C*D*A*B"),
    //.LUTG0("(~C*~(A*~((~B*~D))*~(1)+A*(~B*~D)*~(1)+~(A)*(~B*~D)*1+A*(~B*~D)*1))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000010100000101),
    .INIT_LUTF1(16'b1100010001000100),
    .INIT_LUTG0(16'b0000111100001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2340|_al_u2339  (
    .a({_al_u2339_o,\picorv32_core/mem_rdata_latched [4]}),
    .b({_al_u1536_o,_al_u1483_o_placeOpt_2}),
    .c({_al_u2271_o,_al_u1481_o_placeOpt_2}),
    .d({_al_u1653_o,_al_u2337_o}),
    .e({_al_u2338_o,_al_u1485_o_placeOpt_3}),
    .f({_al_u2340_o,_al_u2339_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~A*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))"),
    //.LUTF1("(~D*~(~0*A*B*C))"),
    //.LUTG0("(~1*~A*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))"),
    //.LUTG1("(~D*~(~1*A*B*C))"),
    .INIT_LUTF0(16'b0100000001010001),
    .INIT_LUTF1(16'b0000000001111111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2342|_al_u2341  (
    .a({\picorv32_core/mem_rdata_latched$1$_placeOpt_1 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_1 }),
    .b({\picorv32_core/mem_rdata_latched [4],_al_u2291_o}),
    .c({_al_u2278_o,\picorv32_core/mem_rdata_latched [6]}),
    .d({_al_u2341_o,_al_u2337_o}),
    .e({\picorv32_core/mem_rdata_latched$0$_placeOpt_4 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .f({_al_u2342_o,_al_u2341_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A)*~((B*C))+D*A*~((B*C))+~(D)*A*(B*C)+D*A*(B*C))"),
    //.LUT1("~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111110000000),
    .INIT_LUT1(16'b0010001001110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2344|picorv32_core/reg6_b20  (
    .a({\picorv32_core/mem_xfer ,\picorv32_core/mem_rdata_latched [31]}),
    .b({\picorv32_core/mem_rdata_latched [31],\picorv32_core/mem_rdata_latched [0]}),
    .c({open_n15662,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [31],\picorv32_core/mem_rdata_latched [12]}),
    .f({_al_u2344_o,open_n15676}),
    .q({open_n15680,\picorv32_core/decoded_imm_uj [20]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B*D)"),
    //.LUT1("(C*~(A*~(~D*~B)))"),
    .INIT_LUT0(16'b0001000100000000),
    .INIT_LUT1(16'b0101000001110000),
    .MODE("LOGIC"))
    \_al_u2345|_al_u2444  (
    .a({_al_u2344_o,_al_u1485_o}),
    .b({_al_u1444_o,_al_u1481_o_placeOpt_4}),
    .c({_al_u1464_o,open_n15681}),
    .d({_al_u1485_o,_al_u1464_o}),
    .f({_al_u2345_o,_al_u2444_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(~(C)*B*~(D)*~(0)+~(C)*~(B)*~(D)*0+C*~(B)*~(D)*0+~(C)*B*~(D)*0+C*B*~(D)*0+~(C)*~(B)*D*0+~(C)*B*D*0))"),
    //.LUT1("(~A*(~(C)*B*~(D)*~(1)+~(C)*~(B)*~(D)*1+C*~(B)*~(D)*1+~(C)*B*~(D)*1+C*B*~(D)*1+~(C)*~(B)*D*1+~(C)*B*D*1))"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000010101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2346 (
    .a({_al_u2344_o,_al_u2344_o}),
    .b({_al_u1481_o_placeOpt_4,_al_u1481_o_placeOpt_4}),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_4 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .d({_al_u1483_o_placeOpt_2,_al_u1483_o_placeOpt_2}),
    .mi({open_n15714,_al_u1485_o_placeOpt_3}),
    .fx({open_n15719,_al_u2346_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A*~B)"),
    //.LUT1("(~A*~(~C*~B))"),
    .INIT_LUT0(16'b0000000100000001),
    .INIT_LUT1(16'b0101010001010100),
    .MODE("LOGIC"))
    \_al_u2347|_al_u2329  (
    .a({_al_u1483_o_placeOpt_1,_al_u1483_o_placeOpt_1}),
    .b({_al_u1481_o_placeOpt_3,_al_u1481_o_placeOpt_3}),
    .c({_al_u1485_o_placeOpt_2,_al_u1485_o_placeOpt_2}),
    .f({_al_u2347_o,_al_u2329_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*D))"),
    //.LUT1("(A*D)"),
    .INIT_LUT0(16'b0100010011001100),
    .INIT_LUT1(16'b1010101000000000),
    .MODE("LOGIC"))
    \_al_u2348|_al_u2367  (
    .a({\picorv32_core/mem_rdata_latched$0$_placeOpt_4 ,_al_u1483_o_placeOpt_2}),
    .b({open_n15744,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .d({\picorv32_core/mem_rdata_latched [12],\picorv32_core/mem_rdata_latched [12]}),
    .f({_al_u2348_o,_al_u2367_o}));
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D)*~(C)*~((A*~B))*~(0)+D*~(C)*~((A*~B))*~(0)+~(D)*C*~((A*~B))*~(0)+D*C*~((A*~B))*~(0)+~(D)*~(C)*(A*~B)*~(0)+D*~(C)*(A*~B)*~(0)+D*C*(A*~B)*~(0)+D*C*~((A*~B))*0+D*C*(A*~B)*0)"),
    //.LUTF1("(~0*~(~B*~(D*~(C*~A))))"),
    //.LUTG0("(~(D)*~(C)*~((A*~B))*~(1)+D*~(C)*~((A*~B))*~(1)+~(D)*C*~((A*~B))*~(1)+D*C*~((A*~B))*~(1)+~(D)*~(C)*(A*~B)*~(1)+D*~(C)*(A*~B)*~(1)+D*C*(A*~B)*~(1)+D*C*~((A*~B))*1+D*C*(A*~B)*1)"),
    //.LUTG1("(~1*~(~B*~(D*~(C*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111011111),
    .INIT_LUTF1(16'b1110111111001100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2349|picorv32_core/reg0_b31  (
    .a({_al_u2345_o,\picorv32_core/n180 }),
    .b({_al_u2346_o,_al_u2351_o}),
    .c({_al_u2347_o,_al_u1569_o}),
    .clk(clk_pad),
    .d({_al_u2348_o,_al_u2349_o}),
    .e({\picorv32_core/mem_rdata_latched [1],_al_u2344_o}),
    .f({_al_u2349_o,open_n15783}),
    .q({open_n15787,\picorv32_core/mem_rdata_q [31]}));  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("B*A*C*~D+B*A*C*D"),
    //.LUTF1("D*~A*~C*B+D*A*~C*B"),
    //.LUTG0("0"),
    //.LUTG1("~D*~A*~C*B+D*~A*~C*B+~D*A*~C*B+D*A*~C*B+~D*~A*C*B+D*~A*C*B+~D*A*C*B+D*A*C*B"),
    .INIT_LUTF0(16'b1000000010000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2350|_al_u1532  (
    .a({open_n15788,\picorv32_core/mem_rdata_latched$0$_placeOpt_2 }),
    .b({\picorv32_core/mem_rdata_latched$1$_placeOpt_3 ,_al_u1481_o}),
    .c({_al_u1483_o_placeOpt_3,_al_u1483_o_placeOpt_3}),
    .d({_al_u1481_o,open_n15791}),
    .e({_al_u1485_o_placeOpt_1,\picorv32_core/mem_rdata_latched$1$_placeOpt_3 }),
    .f({_al_u2350_o,_al_u1532_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~(D*B*A)))"),
    //.LUT1("(D*~(~1*~(A*B*C)))"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2351 (
    .a({\picorv32_core/mem_rdata_latched [12],_al_u1605_o}),
    .b({_al_u1654_o,_al_u1654_o}),
    .c({_al_u1605_o,_al_u2350_o}),
    .d({_al_u2350_o,\picorv32_core/mem_rdata_latched [12]}),
    .mi({open_n15824,_al_u1485_o}),
    .fx({open_n15829,_al_u2351_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A)*~((B*C))+D*A*~((B*C))+~(D)*A*(B*C)+D*A*(B*C))"),
    //.LUT1("~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111110000000),
    .INIT_LUT1(16'b0000111101010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2354|picorv32_core/reg6_b10  (
    .a({\picorv32_core/mem_rdata_q [30],\picorv32_core/mem_rdata_latched [30]}),
    .b({open_n15832,\picorv32_core/mem_rdata_latched$0$_placeOpt_2 }),
    .c({\picorv32_core/mem_rdata_latched [30],\picorv32_core/mem_rdata_latched$1$_placeOpt_3 }),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_xfer_placeOpt_2 ,\picorv32_core/mux79_b1/B0_3 }),
    .f({_al_u2354_o,open_n15846}),
    .q({open_n15850,\picorv32_core/decoded_imm_uj [10]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D)*~(B)*~(C)*~(A)*~(0)+D*~(B)*~(C)*~(A)*~(0)+~(D)*B*~(C)*~(A)*~(0)+D*B*~(C)*~(A)*~(0)+~(D)*~(B)*C*~(A)*~(0)+D*~(B)*C*~(A)*~(0)+~(D)*B*C*~(A)*~(0)+D*B*C*~(A)*~(0)+~(D)*~(B)*~(C)*~(A)*0+D*~(B)*~(C)*~(A)*0+~(D)*B*~(C)*~(A)*0+D*B*~(C)*~(A)*0+~(D)*~(B)*~(C)*A*0+~(D)*B*~(C)*A*0+~(D)*B*C*A*0+D*B*C*A*0)"),
    //.LUT1("(~(D)*~(A)*~(C)*~(B)*~(1)+D*~(A)*~(C)*~(B)*~(1)+~(D)*A*~(C)*~(B)*~(1)+D*A*~(C)*~(B)*~(1)+~(D)*~(A)*C*~(B)*~(1)+D*~(A)*C*~(B)*~(1)+~(D)*A*C*~(B)*~(1)+D*A*C*~(B)*~(1)+~(D)*~(A)*~(C)*~(B)*1+D*~(A)*~(C)*~(B)*1+~(D)*A*~(C)*~(B)*1+D*A*~(C)*~(B)*1+~(D)*~(A)*~(C)*B*1+~(D)*A*~(C)*B*1+~(D)*A*C*B*1+D*A*C*B*1)"),
    .INIT_LUT0(16'b0101010101010101),
    .INIT_LUT1(16'b1000001110001111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2355 (
    .a({_al_u2354_o,_al_u1444_o}),
    .b({_al_u1444_o,_al_u2354_o}),
    .c({\picorv32_core/mem_rdata_latched [12],\picorv32_core/mem_rdata_latched [12]}),
    .d({_al_u1498_o,_al_u1498_o}),
    .mi({open_n15863,_al_u1464_o}),
    .fx({open_n15868,_al_u2355_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*C*~(~A*~(D*~B)))"),
    //.LUTF1("0"),
    //.LUTG0("(1*C*~(~A*~(D*~B)))"),
    //.LUTG1("~D*~A*~B*~C+D*~A*~B*~C+D*A*~B*~C+D*~A*B*~C+D*A*B*~C+~D*~A*~B*C+D*~A*~B*C+D*A*~B*C+D*~A*B*C+D*A*B*C"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1011000010100000),
    .INIT_LUTG1(16'b1111111100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2356|_al_u2357  (
    .a({_al_u1481_o,_al_u2356_o}),
    .b({_al_u1485_o_placeOpt_1,_al_u2355_o}),
    .c({open_n15871,_al_u2273_o}),
    .d({_al_u1483_o_placeOpt_3,\picorv32_core/n98_lutinv }),
    .e({\picorv32_core/mem_rdata_latched [12],\picorv32_core/mem_rdata_latched$0$_placeOpt_2 }),
    .f({_al_u2356_o,_al_u2357_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~D*~C+~A*B*~D*~C+~A*~B*D*~C+~A*B*D*~C+~A*~B*~D*C+~A*B*~D*C+~A*~B*D*C+~A*B*D*C"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("~A*~B*~D*C+~A*B*~D*C+~A*~B*D*C+~A*B*D*C"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0101010101010101),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0101000001010000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2359|_al_u2358  (
    .a({open_n15894,_al_u1485_o_placeOpt_1}),
    .c({_al_u1650_o,_al_u1483_o_placeOpt_3}),
    .d({_al_u2358_o,open_n15899}),
    .e({open_n15900,_al_u1481_o_placeOpt_1}),
    .f({_al_u2359_o,_al_u2358_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*C*D+A*B*C*D"),
    //.LUTF1("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0001110100011101),
    .INIT_LUTG0(16'b1111001111111111),
    .INIT_LUTG1(16'b0001110100011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2363|picorv32_core/reg6_b9  (
    .a({\picorv32_core/mem_rdata_q [29],open_n15921}),
    .b({\picorv32_core/mem_xfer ,\picorv32_core/mem_rdata_latched [0]}),
    .c({\picorv32_core/mem_rdata_latched [29],\picorv32_core/mem_rdata_latched [29]}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({open_n15922,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .e({open_n15923,_al_u1444_o}),
    .f({_al_u2363_o,open_n15939}),
    .q({open_n15943,\picorv32_core/decoded_imm_uj [9]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(~A*~(~B*C)))"),
    //.LUT1("(D*~(C)*~(B)*~(A)+~(D)*~(C)*B*~(A)+D*~(C)*B*~(A)+~(D)*C*B*~(A)+~(D)*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111101000101),
    .INIT_LUT1(16'b0000010111000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2364|picorv32_core/reg0_b29  (
    .a({\picorv32_core/mem_rdata_latched$0$_placeOpt_2 ,_al_u2363_o}),
    .b({_al_u2363_o,_al_u2360_o}),
    .c({\picorv32_core/mux79_b3/B1_0 ,_al_u2353_o}),
    .clk(clk_pad),
    .d({_al_u2358_o,_al_u2368_o}),
    .f({_al_u2364_o,open_n15958}),
    .q({open_n15962,\picorv32_core/mem_rdata_q [29]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(0*~D*~B))"),
    //.LUT1("(C*~A*~(1*~D*~B))"),
    .INIT_LUT0(16'b0101000001010000),
    .INIT_LUT1(16'b0101000001000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2368 (
    .a({_al_u2364_o,_al_u2364_o}),
    .b({_al_u2365_o,_al_u2365_o}),
    .c({_al_u2273_o,_al_u2273_o}),
    .d({_al_u2366_o,_al_u2366_o}),
    .mi({open_n15975,_al_u2367_o}),
    .fx({open_n15980,_al_u2368_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*C*A*~D+B*C*A*~D"),
    //.LUTF1("~A*~C*~B*~D+~A*~C*B*~D"),
    //.LUTG0("0"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000010100000),
    .INIT_LUTF1(16'b0000000000000101),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2370|_al_u2467  (
    .a({_al_u1444_o,_al_u1464_o}),
    .c({_al_u1464_o,_al_u1444_o}),
    .d({\picorv32_core/mux79_b0/B0_3 ,\picorv32_core/n68 [0]}),
    .e({\picorv32_core/mux79_b2/B0_3 ,\picorv32_core/mem_rdata_latched [12]}),
    .f({_al_u2370_o,_al_u2467_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~(C*~(B*D))))"),
    //.LUTF1("(~0*~(~B*A*C*D))"),
    //.LUTG0("(A*~(1*~(C*~(B*D))))"),
    //.LUTG1("(~1*~(~B*A*C*D))"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b1101111111111111),
    .INIT_LUTG0(16'b0010000010100000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2371|_al_u2374  (
    .a({\picorv32_core/mem_rdata_latched [12],\picorv32_core/mem_rdata_latched [12]}),
    .b({\picorv32_core/mux79_b1/B0_3 ,\picorv32_core/mux79_b1/B0_3 }),
    .c({_al_u2370_o,_al_u1483_o_placeOpt_3}),
    .d({_al_u1605_o,_al_u2370_o}),
    .e({_al_u1485_o_placeOpt_1,_al_u1485_o_placeOpt_1}),
    .f({_al_u2371_o,_al_u2374_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A)*~((B*C))+D*A*~((B*C))+~(D)*A*(B*C)+D*A*(B*C))"),
    //.LUT1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111110000000),
    .INIT_LUT1(16'b0000001111001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2372|picorv32_core/reg6_b8  (
    .a({open_n16029,\picorv32_core/mem_rdata_latched [28]}),
    .b({\picorv32_core/mem_xfer_placeOpt_2 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_2 }),
    .c({\picorv32_core/mem_rdata_q [28],\picorv32_core/mem_rdata_latched$1$_placeOpt_3 }),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched [28],\picorv32_core/mux79_b2/B0_3 }),
    .f({_al_u2372_o,open_n16043}),
    .q({open_n16047,\picorv32_core/decoded_imm_uj [8]}));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(A*~(~0*~(B*C))))"),
    //.LUTF1("~A*~D*~C*~B+~A*~D*C*~B+~A*~D*~C*B+~A*D*~C*B+~A*~D*C*B"),
    //.LUTG0("(D*~(A*~(~1*~(B*C))))"),
    //.LUTG1("~A*~D*~C*~B+~A*D*~C*~B+~A*~D*C*~B+~A*D*C*~B+~A*~D*~C*B+~A*D*~C*B+~A*~D*C*B+~A*D*C*B"),
    .INIT_LUTF0(16'b0111111100000000),
    .INIT_LUTF1(16'b0000010001010101),
    .INIT_LUTG0(16'b0101010100000000),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2373|_al_u2353  (
    .a({_al_u2372_o,_al_u2350_o}),
    .b({_al_u2350_o,_al_u1605_o}),
    .c({_al_u2371_o,_al_u1635_o}),
    .d({_al_u1569_o,_al_u1569_o}),
    .e({_al_u2360_o,_al_u1485_o_placeOpt_1}),
    .f({_al_u2373_o,_al_u2353_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(~B*~(D*A))"),
    //.LUTG0("~C*D*A*~B+C*D*A*~B+~C*D*A*B+C*D*A*B"),
    //.LUTG1("(~B*~(D*A))"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000100110011),
    .INIT_LUTG0(16'b1010101000000000),
    .INIT_LUTG1(16'b0001000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2376|_al_u2375  (
    .a({_al_u1579_o,_al_u1485_o_placeOpt_1}),
    .b({_al_u2374_o,open_n16070}),
    .d({_al_u2375_o,_al_u1483_o_placeOpt_3}),
    .e({open_n16075,\picorv32_core/mem_rdata_latched [4]}),
    .f({_al_u2376_o,_al_u2375_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*B*D*~(A*~C))"),
    //.LUTF1("(0*A*D*~(B*C))"),
    //.LUTG0("(1*B*D*~(A*~C))"),
    //.LUTG1("(1*A*D*~(B*C))"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1100010000000000),
    .INIT_LUTG1(16'b0010101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2377|_al_u2410  (
    .a({\picorv32_core/mem_rdata_latched [12],_al_u1444_o}),
    .b({_al_u1444_o,\picorv32_core/mem_rdata_latched [12]}),
    .c({_al_u2372_o,\picorv32_core/n42 [26]}),
    .d({\picorv32_core/n98_lutinv ,\picorv32_core/n98_lutinv }),
    .e({_al_u1464_o,_al_u1464_o}),
    .f({_al_u2377_o,_al_u2410_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTF1("A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("0"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2379|_al_u2430  (
    .a({_al_u2291_o,open_n16118}),
    .c({open_n16121,_al_u1485_o}),
    .d({\picorv32_core/mux79_b2/B0_3 ,\picorv32_core/mux79_b2/B0_3 }),
    .e({_al_u1483_o,_al_u1483_o}),
    .f({_al_u2379_o,_al_u2430_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~0*~C*~(~A*~B)))"),
    //.LUT1("(D*~(~1*~C*~(~A*~B)))"),
    .INIT_LUT0(16'b1111000100000000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2380 (
    .a({_al_u2372_o,_al_u2372_o}),
    .b({_al_u2358_o,_al_u2358_o}),
    .c({_al_u2379_o,_al_u2379_o}),
    .d({_al_u2273_o,_al_u2273_o}),
    .mi({open_n16156,\picorv32_core/mem_rdata_latched$0$_placeOpt_1 }),
    .fx({open_n16161,_al_u2380_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~B*A*C*D)"),
    //.LUT1("(~1*~B*A*C*D)"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2382 (
    .a({\picorv32_core/mux79_b1/B0_3 ,\picorv32_core/mux79_b1/B0_3 }),
    .b({\picorv32_core/mux79_b2/B0_3 ,\picorv32_core/mux79_b2/B0_3 }),
    .c({_al_u1634_o,_al_u1634_o}),
    .d({_al_u2323_o,_al_u2323_o}),
    .mi({open_n16176,\picorv32_core/mux79_b0/B0_3 }),
    .fx({open_n16181,_al_u2382_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~((A*D))+B*C*~((A*D))+~(B)*C*(A*D)+B*C*(A*D))"),
    //.LUT1("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110010011001100),
    .INIT_LUT1(16'b0011010100110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2383|picorv32_core/reg6_b5  (
    .a({\picorv32_core/mem_rdata_q [25],\picorv32_core/mem_rdata_latched [0]}),
    .b({\picorv32_core/mem_rdata_latched [25],\picorv32_core/mem_rdata_latched [2]}),
    .c({\picorv32_core/mem_xfer ,\picorv32_core/mem_rdata_latched [25]}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({open_n16184,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .f({_al_u2383_o,open_n16198}),
    .q({open_n16202,\picorv32_core/decoded_imm_uj [5]}));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~B*~C*~(0*D)))"),
    //.LUTF1("0"),
    //.LUTG0("(A*~(~B*~C*~(1*D)))"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D"),
    .INIT_LUTF0(16'b1010100010101000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0011001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2384|_al_u2385  (
    .a({open_n16203,_al_u2293_o}),
    .b({_al_u2383_o,_al_u2384_o}),
    .c({open_n16204,_al_u2374_o}),
    .d({open_n16207,_al_u2382_o}),
    .e({\picorv32_core/mux81_sel_is_1_o ,\picorv32_core/mem_rdata_latched [2]}),
    .f({_al_u2384_o,_al_u2385_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D*~(~A*~B)))"),
    //.LUT1("(~(B*D)*~(A)*~(C)+~(B*D)*A*~(C)+~(~(B*D))*A*C+~(B*D)*A*C)"),
    .INIT_LUT0(16'b0001000011110000),
    .INIT_LUT1(16'b1010001110101111),
    .MODE("LOGIC"))
    \_al_u2386|_al_u2393  (
    .a({_al_u2383_o,\picorv32_core/mem_do_rinst }),
    .b({_al_u1483_o_placeOpt_3,\picorv32_core/mem_do_prefetch }),
    .c({_al_u1485_o_placeOpt_1,_al_u2383_o}),
    .d({\picorv32_core/mem_rdata_latched [12],_al_u1546_o}),
    .f({_al_u2386_o,_al_u2393_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~0*C*D)))"),
    //.LUT1("(A*~(B*~(~1*C*D)))"),
    .INIT_LUT0(16'b1010001000100010),
    .INIT_LUT1(16'b0010001000100010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2387 (
    .a({_al_u1606_o,_al_u1606_o}),
    .b({_al_u2386_o,_al_u2386_o}),
    .c({_al_u1635_o,_al_u1635_o}),
    .d({_al_u2277_o,_al_u2277_o}),
    .mi({open_n16260,_al_u2383_o}),
    .fx({open_n16265,_al_u2387_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~((~0*~(~B*A)))+~(D)*C*~((~0*~(~B*A)))+~(D)*~(C)*(~0*~(~B*A))+D*~(C)*(~0*~(~B*A))+~(D)*C*(~0*~(~B*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(D*~(C)*~((~1*~(~B*A)))+~(D)*C*~((~1*~(~B*A)))+~(D)*~(C)*(~1*~(~B*A))+D*~(C)*(~1*~(~B*A))+~(D)*C*(~1*~(~B*A)))"),
    //.LUTG1("A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    .INIT_LUTF0(16'b0000111111111101),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000111111110000),
    .INIT_LUTG1(16'b0000111000001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2390|_al_u2389  (
    .a({_al_u2389_o,_al_u1481_o_placeOpt_1}),
    .b({_al_u2383_o,_al_u1483_o_placeOpt_1}),
    .c({_al_u2388_o,\picorv32_core/mem_rdata_latched$0$_placeOpt_1 }),
    .d({open_n16270,\picorv32_core/mem_rdata_latched$1$_placeOpt_1 }),
    .e({_al_u1569_o,_al_u1485_o_placeOpt_2}),
    .f({_al_u2390_o,_al_u2389_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*(~D*~(C)*~(0)+~D*C*~(0)+~(~D)*C*0+~D*C*0))"),
    //.LUTF1("(~(C)*~(B)*~((A*D))*~(0)+C*~(B)*~((A*D))*~(0)+~(C)*B*~((A*D))*~(0)+C*B*~((A*D))*~(0)+C*B*(A*D)*~(0)+C*~(B)*~((A*D))*0+C*B*~((A*D))*0+C*~(B)*(A*D)*0+C*B*(A*D)*0)"),
    //.LUTG0("(B*A*(~D*~(C)*~(1)+~D*C*~(1)+~(~D)*C*1+~D*C*1))"),
    //.LUTG1("(~(C)*~(B)*~((A*D))*~(1)+C*~(B)*~((A*D))*~(1)+~(C)*B*~((A*D))*~(1)+C*B*~((A*D))*~(1)+C*B*(A*D)*~(1)+C*~(B)*~((A*D))*1+C*B*~((A*D))*1+C*~(B)*(A*D)*1+C*B*(A*D)*1)"),
    .INIT_LUTF0(16'b0000000010001000),
    .INIT_LUTF1(16'b1101010111111111),
    .INIT_LUTG0(16'b1000000010000000),
    .INIT_LUTG1(16'b1111000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2391|_al_u2392  (
    .a({_al_u1464_o,_al_u1536_o}),
    .b({_al_u1444_o,_al_u1481_o_placeOpt_1}),
    .c({_al_u2383_o,\picorv32_core/mem_rdata_latched [2]}),
    .d({\picorv32_core/mem_rdata_latched [12],_al_u2391_o}),
    .e({_al_u1485_o_placeOpt_1,_al_u1483_o_placeOpt_3}),
    .f({_al_u2391_o,_al_u2392_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTF1("(~A*~B)"),
    //.LUTG0("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG1("(~A*~B)"),
    .INIT_LUTF0(16'b0011001100110011),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b0001000100010001),
    .INIT_LUTG1(16'b0001000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2395|_al_u2413  (
    .a({_al_u1485_o_placeOpt_2,_al_u1485_o_placeOpt_2}),
    .b({_al_u1481_o_placeOpt_3,_al_u1481_o_placeOpt_3}),
    .e({open_n16319,\picorv32_core/n42 [26]}),
    .f({_al_u2395_o,_al_u2413_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*D*(0*~(B)*~(C)+0*B*~(C)+~(0)*B*C+0*B*C))"),
    //.LUTF1("(A*~B*~D)"),
    //.LUTG0("(A*D*(1*~(B)*~(C)+1*B*~(C)+~(1)*B*C+1*B*C))"),
    //.LUTG1("(A*~B*~D)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000000000100010),
    .INIT_LUTG0(16'b1000101000000000),
    .INIT_LUTG1(16'b0000000000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2396|_al_u2399  (
    .a({_al_u1606_o,_al_u1606_o}),
    .b({_al_u1597_o,\picorv32_core/mem_rdata_latched [3]}),
    .c({open_n16340,_al_u2395_o}),
    .d({_al_u2395_o,_al_u1597_o}),
    .e({open_n16343,\picorv32_core/mux79_b1/B0_3 }),
    .f({_al_u2396_o,_al_u2399_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("C*B*~A*D+C*B*A*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTG0("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0011001111111111),
    .INIT_LUTG0(16'b1111111100111111),
    .INIT_LUTG1(16'b0000000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2397|picorv32_core/reg6_b7  (
    .b({\picorv32_core/mem_xfer ,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .c({open_n16366,\picorv32_core/mem_rdata_latched [0]}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched [27],\picorv32_core/mem_rdata_latched [27]}),
    .e({\picorv32_core/mem_rdata_q [27],\picorv32_core/mem_rdata_latched [6]}),
    .f({_al_u2397_o,open_n16382}),
    .q({open_n16386,\picorv32_core/decoded_imm_uj [7]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~(A*C*~(B*~D)))"),
    //.LUT1("(~1*~(A*C*~(B*~D)))"),
    .INIT_LUT0(16'b0101111111011111),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2398 (
    .a({_al_u2389_o,_al_u2389_o}),
    .b({_al_u2396_o,_al_u2396_o}),
    .c({_al_u1569_o,_al_u1569_o}),
    .d({_al_u2371_o,_al_u2371_o}),
    .mi({open_n16399,_al_u2397_o}),
    .fx({open_n16404,_al_u2398_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~A*~(C*~(~0*~B))))"),
    //.LUTF1("(A*~(~C*~(D*~(~0*~B))))"),
    //.LUTG0("(D*~(~A*~(C*~(~1*~B))))"),
    //.LUTG1("(A*~(~C*~(D*~(~1*~B))))"),
    .INIT_LUTF0(16'b1110101000000000),
    .INIT_LUTF1(16'b1010100010100000),
    .INIT_LUTG0(16'b1111101000000000),
    .INIT_LUTG1(16'b1010101010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2400|_al_u1645  (
    .a({\picorv32_core/mux79_b1/B0_3 ,_al_u1638_o}),
    .b({_al_u1439_o,_al_u1439_o}),
    .c({_al_u1638_o,_al_u1637_o}),
    .d({_al_u1637_o,\picorv32_core/mem_rdata_latched [2]}),
    .e({_al_u1088_o,_al_u1088_o}),
    .f({_al_u2400_o,\picorv32_core/sel10_b0/B1_1 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C)*~(B)*~(A)*~(D)*~(0)+C*~(B)*~(A)*~(D)*~(0)+~(C)*B*~(A)*~(D)*~(0)+C*B*~(A)*~(D)*~(0)+~(C)*~(B)*A*~(D)*~(0)+C*~(B)*A*~(D)*~(0)+~(C)*B*A*~(D)*~(0)+C*B*A*~(D)*~(0)+C*~(B)*~(A)*D*~(0)+~(C)*B*~(A)*D*~(0)+~(C)*~(B)*A*D*~(0)+C*~(B)*A*D*~(0)+~(C)*B*A*D*~(0)+~(C)*~(B)*~(A)*~(D)*0+C*~(B)*~(A)*~(D)*0+~(C)*B*~(A)*~(D)*0+~(C)*~(B)*A*~(D)*0+C*~(B)*A*~(D)*0+~(C)*B*A*~(D)*0+C*~(B)*~(A)*D*0+~(C)*B*~(A)*D*0+~(C)*~(B)*A*D*0+C*~(B)*A*D*0+~(C)*B*A*D*0)"),
    //.LUT1("(~(C)*~(A)*~(B)*~(D)*~(1)+C*~(A)*~(B)*~(D)*~(1)+~(C)*A*~(B)*~(D)*~(1)+C*A*~(B)*~(D)*~(1)+~(C)*~(A)*B*~(D)*~(1)+C*~(A)*B*~(D)*~(1)+~(C)*A*B*~(D)*~(1)+C*A*B*~(D)*~(1)+C*~(A)*~(B)*D*~(1)+~(C)*A*~(B)*D*~(1)+~(C)*~(A)*B*D*~(1)+C*~(A)*B*D*~(1)+~(C)*A*B*D*~(1)+~(C)*~(A)*~(B)*~(D)*1+C*~(A)*~(B)*~(D)*1+~(C)*A*~(B)*~(D)*1+~(C)*~(A)*B*~(D)*1+C*~(A)*B*~(D)*1+~(C)*A*B*~(D)*1+C*~(A)*~(B)*D*1+~(C)*A*~(B)*D*1+~(C)*~(A)*B*D*1+C*~(A)*B*D*1+~(C)*A*B*D*1)"),
    .INIT_LUT0(16'b0011111011111111),
    .INIT_LUT1(16'b0101111001011111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2401 (
    .a({_al_u2400_o,_al_u2397_o}),
    .b({_al_u2397_o,_al_u2400_o}),
    .c({_al_u1650_o,_al_u1650_o}),
    .d({\picorv32_core/mux81_sel_is_1_o ,\picorv32_core/mux81_sel_is_1_o }),
    .mi({open_n16441,_al_u2329_o}),
    .fx({open_n16446,_al_u2401_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(0*C*D*~(A*B))"),
    //.LUT1("(1*C*D*~(B*A))"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0111000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2402 (
    .a({_al_u2397_o,_al_u1444_o}),
    .b({_al_u1444_o,_al_u2397_o}),
    .c({\picorv32_core/mem_rdata_latched [12],\picorv32_core/mem_rdata_latched [12]}),
    .d({\picorv32_core/n98_lutinv ,\picorv32_core/n98_lutinv }),
    .mi({open_n16461,_al_u1464_o}),
    .fx({open_n16466,_al_u2402_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~A*~(0*~(~B*~C)))"),
    //.LUT1("(D*~A*~(1*~(~B*~C)))"),
    .INIT_LUT0(16'b0101010100000000),
    .INIT_LUT1(16'b0000000100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2404 (
    .a({_al_u2399_o,_al_u2399_o}),
    .b({_al_u2403_o,_al_u2403_o}),
    .c({_al_u2402_o,_al_u2402_o}),
    .d({_al_u2401_o,_al_u2401_o}),
    .mi({open_n16481,_al_u1536_o}),
    .fx({open_n16486,_al_u2404_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*A)"),
    //.LUT1("(D*A)"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010101000000000),
    .MODE("LOGIC"))
    \_al_u2405|_al_u2323  (
    .a({_al_u2323_o,_al_u1483_o_placeOpt_1}),
    .b({open_n16489,_al_u1485_o_placeOpt_2}),
    .d({\picorv32_core/mem_rdata_latched [3],open_n16494}),
    .f({_al_u2405_o,_al_u2323_o}));
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*B*~C*~A+D*B*~C*~A+D*B*C*~A+~D*B*~C*A+D*B*~C*A+D*B*C*A"),
    //.LUTF1("A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG1("A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110000001100),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b1111111111111111),
    .INIT_LUTG1(16'b1010101010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2406|picorv32_core/reg0_b27  (
    .a({_al_u2293_o,open_n16513}),
    .b({open_n16514,_al_u1569_o}),
    .c({_al_u1579_o,_al_u2404_o}),
    .clk(clk_pad),
    .d({_al_u2374_o,_al_u2406_o}),
    .e({_al_u2405_o,_al_u2398_o}),
    .f({_al_u2406_o,open_n16531}),
    .q({open_n16535,\picorv32_core/mem_rdata_q [27]}));  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("~((0*A)*~((B*D))*~(C)+(0*A)*(B*D)*~(C)+~((0*A))*(B*D)*C+(0*A)*(B*D)*C)"),
    //.LUTF1("(B*~(A*~D*~(~0*~C)))"),
    //.LUTG0("~((1*A)*~((B*D))*~(C)+(1*A)*(B*D)*~(C)+~((1*A))*(B*D)*C+(1*A)*(B*D)*C)"),
    //.LUTG1("(B*~(A*~D*~(~1*~C)))"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b1100110001001100),
    .INIT_LUTG0(16'b0011010111110101),
    .INIT_LUTG1(16'b1100110001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2412|_al_u2411  (
    .a({_al_u2411_o,\picorv32_core/n42 [26]}),
    .b({_al_u1536_o,_al_u1481_o_placeOpt_3}),
    .c({_al_u2408_o,_al_u1483_o_placeOpt_1}),
    .d({_al_u2410_o,\picorv32_core/mem_rdata_latched [5]}),
    .e({_al_u1481_o_placeOpt_3,_al_u1485_o_placeOpt_2}),
    .f({_al_u2412_o,_al_u2411_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*C*~D)"),
    //.LUT1("(A*~(C*~(B*D)))"),
    .INIT_LUT0(16'b0000000010100000),
    .INIT_LUT1(16'b1000101000001010),
    .MODE("LOGIC"))
    \_al_u2414|_al_u1593  (
    .a({_al_u1606_o,\picorv32_core/mem_rdata_latched$0$_placeOpt_1 }),
    .b({\picorv32_core/mem_rdata_latched [2],open_n16558}),
    .c({_al_u2413_o,\picorv32_core/mem_rdata_latched$1$_placeOpt_1 }),
    .d({_al_u1597_o,\picorv32_core/mem_rdata_latched [2]}),
    .f({_al_u2414_o,_al_u1593_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*(D*~(A)*~(0)+D*A*~(0)+~(D)*A*0+D*A*0)))"),
    //.LUT1("(B*~(C*(D*~(A)*~(1)+D*A*~(1)+~(D)*A*1+D*A*1)))"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b0100110001001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2415 (
    .a({\picorv32_core/n42 [26],\picorv32_core/n42 [26]}),
    .b({_al_u1481_o_placeOpt_3,_al_u1481_o_placeOpt_3}),
    .c({_al_u1483_o_placeOpt_1,_al_u1483_o_placeOpt_1}),
    .d({\picorv32_core/mux79_b0/B0_3 ,\picorv32_core/mux79_b0/B0_3 }),
    .mi({open_n16591,_al_u1485_o_placeOpt_2}),
    .fx({open_n16596,_al_u2415_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(~0*A*~D)))"),
    //.LUT1("(C*~(B*~(~1*A*~D)))"),
    .INIT_LUT0(16'b0011000010110000),
    .INIT_LUT1(16'b0011000000110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2416 (
    .a({\picorv32_core/n42 [26],\picorv32_core/n42 [26]}),
    .b({_al_u2415_o,_al_u2415_o}),
    .c({_al_u2414_o,_al_u2414_o}),
    .d({_al_u2371_o,_al_u2371_o}),
    .mi({open_n16611,_al_u1483_o_placeOpt_1}),
    .fx({open_n16616,_al_u2416_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*((~A*D)*~(C)*~(B)+(~A*D)*C*~(B)+~((~A*D))*C*B+(~A*D)*C*B))"),
    //.LUT1("(~1*((~B*D)*~(A)*~(C)+(~B*D)*A*~(C)+~((~B*D))*A*C+(~B*D)*A*C))"),
    .INIT_LUT0(16'b1101000111000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2417 (
    .a({\picorv32_core/mem_rdata_latched [5],_al_u1481_o_placeOpt_3}),
    .b({_al_u1481_o_placeOpt_3,_al_u1483_o_placeOpt_1}),
    .c({_al_u1483_o_placeOpt_1,\picorv32_core/mem_rdata_latched [5]}),
    .d({\picorv32_core/mux79_b0/B0_3 ,\picorv32_core/mux79_b0/B0_3 }),
    .mi({open_n16631,_al_u1485_o_placeOpt_2}),
    .fx({open_n16636,_al_u2417_o}));
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~0*~A)*~(D*~C*~B))"),
    //.LUTF1("(D*~(C*A)*~(0*~B))"),
    //.LUTG0("(~(~1*~A)*~(D*~C*~B))"),
    //.LUTG1("(D*~(C*A)*~(1*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100010101010),
    .INIT_LUTF1(16'b0101111100000000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b0100110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2418|picorv32_core/reg0_b26  (
    .a({_al_u2417_o,_al_u1569_o}),
    .b({_al_u2389_o,_al_u2412_o}),
    .c({_al_u1650_o,_al_u2416_o}),
    .clk(clk_pad),
    .d({_al_u1569_o,_al_u2418_o}),
    .e({\picorv32_core/n42 [26],\picorv32_core/n42 [26]}),
    .f({_al_u2418_o,open_n16655}),
    .q({open_n16659,\picorv32_core/mem_rdata_q [26]}));  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D"),
    //.LUTF1("~A*~B*~C*D+~A*B*~C*D"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D"),
    //.LUTG1("~A*~B*~C*D+~A*B*~C*D"),
    .INIT_LUTF0(16'b0000000000001010),
    .INIT_LUTF1(16'b0000010100000000),
    .INIT_LUTG0(16'b0000000000001010),
    .INIT_LUTG1(16'b0000010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2420|_al_u2366  (
    .a({\picorv32_core/mem_rdata_latched [12],\picorv32_core/mem_rdata_latched [12]}),
    .c({_al_u1605_o,_al_u1485_o}),
    .d({_al_u1481_o_placeOpt_4,_al_u1481_o_placeOpt_4}),
    .f({_al_u2420_o,_al_u2366_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~A*~C*B+D*~A*~C*B+~D*A*~C*B+D*A*~C*B+~D*~A*C*B+D*~A*C*B"),
    //.LUTF1("(D*~B)"),
    //.LUTG0("~D*A*C*~B+D*A*C*~B+~D*~A*~C*B+D*~A*~C*B+~D*A*~C*B+D*A*~C*B+~D*~A*C*B+D*~A*C*B+~D*A*C*B+D*A*C*B"),
    //.LUTG1("(D*~B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100110001001100),
    .INIT_LUTF1(16'b0011001100000000),
    .INIT_LUTG0(16'b1110110011101100),
    .INIT_LUTG1(16'b0011001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2421|picorv32_core/reg6_b19  (
    .a({open_n16686,\picorv32_core/mem_rdata_latched [0]}),
    .b({\picorv32_core/n180 ,\picorv32_core/mem_rdata_latched [12]}),
    .c({open_n16687,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched [19],open_n16688}),
    .e({open_n16689,\picorv32_core/mem_rdata_latched [19]}),
    .f({_al_u2421_o,open_n16705}),
    .q({open_n16709,\picorv32_core/decoded_imm_uj [19]}));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("A*~B*C*~D+A*B*C*~D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("~B*D*~C*A+B*D*~C*A+~B*D*C*A+B*D*C*A"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010000010100000),
    .INIT_LUTG0(16'b1010101000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2424|_al_u2365  (
    .a({\picorv32_core/n98_lutinv ,\picorv32_core/n98_lutinv }),
    .c({_al_u1536_o,open_n16712}),
    .d({open_n16715,_al_u1464_o}),
    .e({_al_u2295_o,\picorv32_core/mem_rdata_latched [12]}),
    .f({_al_u2424_o,_al_u2365_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~D*~(0*B*~C))"),
    //.LUTF1("0"),
    //.LUTG0("(~A*~D*~(1*B*~C))"),
    //.LUTG1("C*A*~D*~B+~C*~A*D*~B+~C*A*D*~B+C*A*D*~B+C*A*~D*B+~C*~A*D*B+~C*A*D*B+C*A*D*B"),
    .INIT_LUTF0(16'b0000000001010101),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000001010001),
    .INIT_LUTG1(16'b1010111110100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2425|_al_u2426  (
    .a({_al_u1483_o_placeOpt_3,_al_u2425_o}),
    .b({open_n16736,\picorv32_core/mux79_b3/B1_0 }),
    .c({_al_u1481_o,_al_u2420_o}),
    .d({\picorv32_core/mux79_b3/B1_0 ,_al_u2424_o}),
    .e({_al_u1536_o,_al_u1606_o}),
    .f({_al_u2425_o,_al_u2426_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B)"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~B)"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000001100000011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000011),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2427|_al_u2270  (
    .b({_al_u1597_o,\picorv32_core/mux79_b0/B0_3 }),
    .c({open_n16761,\picorv32_core/mux79_b2/B0_3 }),
    .e({_al_u1650_o,open_n16766}),
    .f({_al_u2427_o,_al_u2270_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(~(D)*~(B)*~(C)*~(0)+D*~(B)*~(C)*~(0)+~(D)*B*~(C)*~(0)+~(D)*B*C*~(0)+D*B*C*~(0)+~(D)*B*C*0+D*B*C*0))"),
    //.LUTF1("~((B*A*~D)*~(C)*~(0)+(B*A*~D)*C*~(0)+~((B*A*~D))*C*0+(B*A*~D)*C*0)"),
    //.LUTG0("(A*(~(D)*~(B)*~(C)*~(1)+D*~(B)*~(C)*~(1)+~(D)*B*~(C)*~(1)+~(D)*B*C*~(1)+D*B*C*~(1)+~(D)*B*C*1+D*B*C*1))"),
    //.LUTG1("~((B*A*~D)*~(C)*~(1)+(B*A*~D)*C*~(1)+~((B*A*~D))*C*1+(B*A*~D)*C*1)"),
    .INIT_LUTF0(16'b1000001010001010),
    .INIT_LUTF1(16'b1111111101110111),
    .INIT_LUTG0(16'b1000000010000000),
    .INIT_LUTG1(16'b0000111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2431|_al_u2429  (
    .a({_al_u2430_o,\picorv32_core/mux79_b2/B0_3 }),
    .b({\picorv32_core/mem_rdata_latched [1],_al_u1481_o_placeOpt_4}),
    .c({_al_u2429_o,_al_u1483_o}),
    .d({_al_u2420_o,_al_u2295_o}),
    .e({\picorv32_core/mem_rdata_latched$0$_placeOpt_4 ,_al_u1485_o}),
    .f({_al_u2431_o,_al_u2429_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*A*(~(D)*~(C)*~(0)+D*~(C)*~(0)+D*C*0))"),
    //.LUT1("(~A*B*(~(C)*~(D)*~(1)+C*~(D)*~(1)+C*D*1))"),
    .INIT_LUT0(16'b0000001000000010),
    .INIT_LUT1(16'b0100000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2433 (
    .a({_al_u1481_o_placeOpt_1,\picorv32_core/mux79_b1/B0_3 }),
    .b({\picorv32_core/mux79_b1/B0_3 ,_al_u1481_o_placeOpt_1}),
    .c({_al_u2370_o,_al_u1483_o_placeOpt_1}),
    .d({_al_u1483_o_placeOpt_1,_al_u2370_o}),
    .mi({open_n16821,_al_u1485_o_placeOpt_2}),
    .fx({open_n16826,_al_u2433_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(~(D)*~(A)*~(C)*~(0)+D*~(A)*~(C)*~(0)+~(D)*A*~(C)*~(0)+~(D)*~(A)*C*~(0)+D*~(A)*C*~(0)+~(D)*~(A)*C*0+D*~(A)*C*0))"),
    //.LUTF1("(A*B*~(~C*~(~0*~D)))"),
    //.LUTG0("(B*(~(D)*~(A)*~(C)*~(1)+D*~(A)*~(C)*~(1)+~(D)*A*~(C)*~(1)+~(D)*~(A)*C*~(1)+D*~(A)*C*~(1)+~(D)*~(A)*C*1+D*~(A)*C*1))"),
    //.LUTG1("(A*B*~(~C*~(~1*~D)))"),
    .INIT_LUTF0(16'b0100010001001100),
    .INIT_LUTF1(16'b1000000010001000),
    .INIT_LUTG0(16'b0100000001000000),
    .INIT_LUTG1(16'b1000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2434|_al_u2454  (
    .a({_al_u1481_o_placeOpt_2,_al_u1481_o_placeOpt_2}),
    .b({\picorv32_core/mux79_b1/B0_3 ,\picorv32_core/mux79_b1/B0_3 }),
    .c({_al_u1483_o_placeOpt_2,_al_u1483_o_placeOpt_2}),
    .d({_al_u2295_o,_al_u2295_o}),
    .e({_al_u1485_o_placeOpt_3,_al_u1485_o_placeOpt_3}),
    .f({_al_u2434_o,_al_u2454_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*A*D*~(~C*B))"),
    //.LUTF1("(~0*C*(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D))"),
    //.LUTG0("(~1*A*D*~(~C*B))"),
    //.LUTG1("(~1*C*(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D))"),
    .INIT_LUTF0(16'b1010001000000000),
    .INIT_LUTF1(16'b1100000001010000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2435|_al_u2388  (
    .a({_al_u1481_o_placeOpt_3,\picorv32_core/mem_rdata_latched [12]}),
    .b({\picorv32_core/mux79_b1/B0_3 ,_al_u1481_o_placeOpt_3}),
    .c({_al_u1650_o,_al_u1483_o_placeOpt_1}),
    .d({_al_u1483_o_placeOpt_1,_al_u1650_o}),
    .e({_al_u1485_o_placeOpt_2,_al_u1485_o_placeOpt_2}),
    .f({_al_u2435_o,_al_u2388_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A)*~((B*C))+D*A*~((B*C))+~(D)*A*(B*C)+D*A*(B*C))"),
    //.LUT1("(D*~B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111110000000),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2436|picorv32_core/reg6_b16  (
    .a({open_n16873,\picorv32_core/mem_rdata_latched [16]}),
    .b({\picorv32_core/n180 ,\picorv32_core/mem_rdata_latched [0]}),
    .c({open_n16874,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched [16],\picorv32_core/mem_rdata_latched [12]}),
    .f({_al_u2436_o,open_n16888}),
    .q({open_n16892,\picorv32_core/decoded_imm_uj [16]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(A*~(~B*~(0*~C))))"),
    //.LUTF1("(~A*~B*~(0*~(~C*~D)))"),
    //.LUTG0("~(D*~(A*~(~B*~(1*~C))))"),
    //.LUTG1("(~A*~B*~(1*~(~C*~D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100011111111),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b1000101011111111),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2437|picorv32_core/reg8_b1  (
    .a({_al_u2436_o,_al_u1606_o}),
    .b({_al_u2435_o,_al_u1597_o}),
    .c({_al_u2434_o,_al_u2420_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u2433_o,_al_u2437_o}),
    .e({_al_u1536_o,_al_u2400_o}),
    .f({_al_u2437_o,open_n16908}),
    .q({open_n16912,\picorv32_core/decoded_rs1 [1]}));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*(~(B)*~(A)*~(0)+B*A*~(0)+B*A*0))"),
    //.LUTF1("(~A*~C*~(0*B*~D))"),
    //.LUTG0("(D*C*(~(B)*~(A)*~(1)+B*A*~(1)+B*A*1))"),
    //.LUTG1("(~A*~C*~(1*B*~D))"),
    .INIT_LUTF0(16'b1001000000000000),
    .INIT_LUTF1(16'b0000010100000101),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000010100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2441|_al_u2440  (
    .a({_al_u2440_o,_al_u1483_o_placeOpt_2}),
    .b({\picorv32_core/mux79_b0/B1_0 ,_al_u1481_o_placeOpt_4}),
    .c({_al_u2297_o,_al_u1536_o}),
    .d({_al_u2420_o,\picorv32_core/mux79_b0/B0_3 }),
    .e({_al_u1606_o,_al_u1485_o}),
    .f({_al_u2441_o,_al_u2440_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(0*~(~B*~(A*~C))))"),
    //.LUTF1("(C*A*~(~B*~(~0*~D)))"),
    //.LUTG0("~(~D*~(1*~(~B*~(A*~C))))"),
    //.LUTG1("(C*A*~(~B*~(~1*~D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b1000000010100000),
    .INIT_LUTG0(16'b1111111111001110),
    .INIT_LUTG1(16'b1000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2443|picorv32_core/reg7_b4  (
    .a({\picorv32_core/mem_rdata_latched [0],_al_u2422_o}),
    .b({\picorv32_core/mem_rdata_latched$1$_placeOpt_4 ,_al_u2444_o}),
    .c({_al_u1464_o,_al_u1605_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mux81_sel_is_1_o ,_al_u2443_o}),
    .e({_al_u1481_o_placeOpt_4,_al_u1606_o}),
    .f({_al_u2443_o,open_n16950}),
    .q({open_n16954,\picorv32_core/decoded_rd [4]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~D*~C*~(0*~B))"),
    //.LUTF1("(A*C*~(~B*~(0*~D)))"),
    //.LUTG0("~(~A*~D*~C*~(1*~B))"),
    //.LUTG1("(A*C*~(~B*~(1*~D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111010),
    .INIT_LUTF1(16'b1000000010000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1000000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2446|picorv32_core/reg7_b3  (
    .a({_al_u1444_o,_al_u2447_o}),
    .b({_al_u2291_o,\picorv32_core/n180 }),
    .c({_al_u1606_o,_al_u2446_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u1605_o,_al_u2424_o}),
    .e({\picorv32_core/n98_lutinv ,_al_u1444_o}),
    .f({_al_u2446_o,open_n16970}),
    .q({open_n16974,\picorv32_core/decoded_rd [3]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(~(D)*A*~(B)*~(0)+D*A*~(B)*~(0)+~(D)*A*~(B)*0+D*A*~(B)*0+D*~(A)*B*0+~(D)*A*B*0+D*A*B*0))"),
    //.LUT1("(~B*(~(D)*C*~(A)*~(1)+D*C*~(A)*~(1)+~(D)*C*~(A)*1+D*C*~(A)*1+D*~(C)*A*1+~(D)*C*A*1+D*C*A*1))"),
    .INIT_LUT0(16'b0000001000000010),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2447 (
    .a({\picorv32_core/mem_rdata_latched$0$_placeOpt_3 ,_al_u2291_o}),
    .b({\picorv32_core/mem_rdata_latched [1],\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }),
    .c({_al_u2291_o,\picorv32_core/mem_rdata_latched [1]}),
    .d({_al_u1625_o,_al_u1625_o}),
    .mi({open_n16987,_al_u1444_o}),
    .fx({open_n16992,_al_u2447_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*C*D*~(0*A))"),
    //.LUTF1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+~A*D*C*~B+~A*D*~C*B+A*D*~C*B+~A*D*C*B"),
    //.LUTG0("(~B*C*D*~(1*A))"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+~A*D*C*~B"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b0101111100010011),
    .INIT_LUTG0(16'b0001000000000000),
    .INIT_LUTG1(16'b0001001100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2449|_al_u2315  (
    .a({\picorv32_core/mux79_b2/B0_3 ,_al_u1654_o}),
    .b({_al_u2430_o,\picorv32_core/mem_rdata_latched [2]}),
    .c({_al_u2291_o,\picorv32_core/n98_lutinv }),
    .d({_al_u1596_o,_al_u1596_o}),
    .e({\picorv32_core/mem_rdata_latched [2],\picorv32_core/mem_rdata_latched [12]}),
    .f({_al_u2449_o,_al_u2315_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(~(D)*~(A)*~(B)*~(0)+D*~(A)*~(B)*~(0)+~(D)*A*~(B)*~(0)+~(D)*~(A)*B*~(0)+D*~(A)*B*~(0)+~(D)*~(A)*B*0+D*~(A)*B*0))"),
    //.LUT1("(A*(~(D)*~(B)*~(C)*~(1)+D*~(B)*~(C)*~(1)+~(D)*B*~(C)*~(1)+~(D)*~(B)*C*~(1)+D*~(B)*C*~(1)+~(D)*~(B)*C*1+D*~(B)*C*1))"),
    .INIT_LUT0(16'b0101000001110000),
    .INIT_LUT1(16'b0010000000100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2450 (
    .a({\picorv32_core/mux79_b2/B0_3 ,_al_u1481_o_placeOpt_2}),
    .b({_al_u1481_o_placeOpt_2,_al_u1483_o_placeOpt_2}),
    .c({_al_u1483_o_placeOpt_2,\picorv32_core/mux79_b2/B0_3 }),
    .d({_al_u2295_o,_al_u2295_o}),
    .mi({open_n17029,_al_u1485_o_placeOpt_3}),
    .fx({open_n17034,_al_u2450_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~((A*D))*~(C)*~(B)*~(0)+~((A*D))*C*~(B)*~(0)+(A*D)*C*~(B)*~(0)+~((A*D))*~(C)*B*~(0)+(A*D)*~(C)*B*~(0)+~((A*D))*C*B*~(0)+(A*D)*C*B*~(0)+~((A*D))*~(C)*~(B)*0+~((A*D))*C*~(B)*0+(A*D)*C*~(B)*0+~((A*D))*~(C)*B*0+(A*D)*~(C)*B*0)"),
    //.LUT1("(~((A*D))*~(C)*~(B)*~(1)+~((A*D))*C*~(B)*~(1)+(A*D)*C*~(B)*~(1)+~((A*D))*~(C)*B*~(1)+(A*D)*~(C)*B*~(1)+~((A*D))*C*B*~(1)+(A*D)*C*B*~(1)+~((A*D))*~(C)*~(B)*1+~((A*D))*C*~(B)*1+(A*D)*C*~(B)*1+~((A*D))*~(C)*B*1+(A*D)*~(C)*B*1)"),
    .INIT_LUT0(16'b1111110111111111),
    .INIT_LUT1(16'b0011110100111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2451 (
    .a({\picorv32_core/mem_rdata_latched [4],\picorv32_core/mem_rdata_latched [4]}),
    .b({\picorv32_core/mem_rdata_latched$0$_placeOpt_4 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .c({\picorv32_core/mem_rdata_latched [1],\picorv32_core/mem_rdata_latched [1]}),
    .d({_al_u2291_o,_al_u2291_o}),
    .mi({open_n17049,\picorv32_core/mux79_b2/B0_3 }),
    .fx({open_n17054,_al_u2451_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(~0*~(~C*D))))"),
    //.LUT1("(B*~(A*~(~1*~(~C*D))))"),
    .INIT_LUT0(16'b1100010011001100),
    .INIT_LUT1(16'b0100010001000100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2453 (
    .a({_al_u1481_o_placeOpt_2,_al_u1481_o_placeOpt_2}),
    .b({_al_u2400_o,_al_u2400_o}),
    .c({\picorv32_core/mem_rdata_latched [2],\picorv32_core/mem_rdata_latched [2]}),
    .d({_al_u1596_o,_al_u1596_o}),
    .mi({open_n17069,_al_u1483_o_placeOpt_2}),
    .fx({open_n17074,_al_u2453_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~((B*D))*~(C)*~(A)*~(0)+~((B*D))*C*~(A)*~(0)+(B*D)*C*~(A)*~(0)+~((B*D))*~(C)*A*~(0)+(B*D)*~(C)*A*~(0)+~((B*D))*C*A*~(0)+(B*D)*C*A*~(0)+~((B*D))*~(C)*~(A)*0+~((B*D))*C*~(A)*0+(B*D)*C*~(A)*0+~((B*D))*~(C)*A*0+(B*D)*~(C)*A*0)"),
    //.LUT1("(~((A*D))*~(C)*~(B)*~(1)+~((A*D))*C*~(B)*~(1)+(A*D)*C*~(B)*~(1)+~((A*D))*~(C)*B*~(1)+(A*D)*~(C)*B*~(1)+~((A*D))*C*B*~(1)+(A*D)*C*B*~(1)+~((A*D))*~(C)*~(B)*1+~((A*D))*C*~(B)*1+(A*D)*C*~(B)*1+~((A*D))*~(C)*B*1+(A*D)*~(C)*B*1)"),
    .INIT_LUT0(16'b1111101111111111),
    .INIT_LUT1(16'b0011110100111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2455 (
    .a({\picorv32_core/mem_rdata_latched [3],\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .b({\picorv32_core/mem_rdata_latched$0$_placeOpt_4 ,\picorv32_core/mem_rdata_latched [3]}),
    .c({\picorv32_core/mem_rdata_latched$1$_placeOpt_1 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_1 }),
    .d({_al_u2291_o,_al_u2291_o}),
    .mi({open_n17089,\picorv32_core/mux79_b1/B0_3 }),
    .fx({open_n17094,_al_u2455_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B*(C*~(A)*~(0)+C*A*~(0)+~(C)*A*0+C*A*0)))"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(D*~(B*(C*~(A)*~(1)+C*A*~(1)+~(C)*A*1+C*A*1)))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1100111111001100),
    .INIT_LUTG0(16'b0111011100000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2461|_al_u2458  (
    .a({open_n17097,_al_u2457_o}),
    .b({\picorv32_core/mem_rdata_latched$1$_placeOpt_3 ,_al_u1602_o}),
    .c({_al_u1483_o_placeOpt_3,_al_u1498_o}),
    .d({_al_u1485_o_placeOpt_1,\picorv32_core/n98_lutinv }),
    .e({_al_u2457_o,\picorv32_core/mem_rdata_latched [12]}),
    .f({_al_u2461_o,_al_u2458_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*~(A*C*B))"),
    //.LUTF1("(C*~(~B*~(~0*~(~A*~D))))"),
    //.LUTG0("(~1*D*~(A*C*B))"),
    //.LUTG1("(C*~(~B*~(~1*~(~A*~D))))"),
    .INIT_LUTF0(16'b0111111100000000),
    .INIT_LUTF1(16'b1111000011100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2462|_al_u2459  (
    .a({_al_u2459_o,\picorv32_core/mux79_b1/B0_3 }),
    .b({_al_u2461_o,_al_u1634_o}),
    .c({_al_u2460_o,_al_u2270_o}),
    .d({_al_u2458_o,_al_u2375_o}),
    .e({\picorv32_core/mem_rdata_latched$1$_placeOpt_3 ,_al_u1481_o}),
    .f({_al_u2462_o,_al_u2459_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~0*~(B*~(A*D))))"),
    //.LUT1("(C*~(~1*~(B*~(A*D))))"),
    .INIT_LUT0(16'b0100000011000000),
    .INIT_LUT1(16'b1111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2464 (
    .a({\picorv32_core/mux79_b1/B0_3 ,\picorv32_core/mux79_b1/B0_3 }),
    .b({\picorv32_core/mem_rdata_latched [2],\picorv32_core/mem_rdata_latched [2]}),
    .c({_al_u2323_o,_al_u2323_o}),
    .d({_al_u2370_o,_al_u2370_o}),
    .mi({open_n17154,_al_u1481_o_placeOpt_1}),
    .fx({open_n17159,_al_u2464_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~(0*~B*~A)))"),
    //.LUTF1("0"),
    //.LUTG0("(D*~(~C*~(1*~B*~A)))"),
    //.LUTG1("D*B*C*~A+D*B*C*A"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000100000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2466|_al_u2468  (
    .a({open_n17162,_al_u2466_o}),
    .b({_al_u1444_o,_al_u2467_o}),
    .c({_al_u2465_o,_al_u2464_o}),
    .d({_al_u1464_o,_al_u2273_o}),
    .e({\picorv32_core/mem_rdata_latched [12],\picorv32_core/n98_lutinv }),
    .f({_al_u2466_o,_al_u2468_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~(~0*~(~A*B)))"),
    //.LUTF1("~D*~A*~C*~B+D*~A*~C*~B+~D*~A*C*~B+D*~A*C*~B"),
    //.LUTG0("(~D*~C*~(~1*~(~A*B)))"),
    //.LUTG1("~D*~A*~C*~B+D*~A*~C*~B+~D*~A*C*~B"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2470|_al_u2469  (
    .a({_al_u2469_o,_al_u1483_o_placeOpt_1}),
    .b({\picorv32_core/mem_rdata_latched$0$_placeOpt_1 ,_al_u1481_o_placeOpt_3}),
    .c({_al_u2329_o,_al_u2465_o}),
    .d({_al_u1569_o,\picorv32_core/mem_rdata_latched$1$_placeOpt_1 }),
    .e({\picorv32_core/mem_rdata_latched$1$_placeOpt_1 ,_al_u1485_o_placeOpt_2}),
    .f({_al_u2470_o,_al_u2469_o}));
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(~0*~A)*~(~C*~(B*~D)))"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*B*C*D"),
    //.LUTG0("~(~(~1*~A)*~(~C*~(B*~D)))"),
    //.LUTG1("A*B*~C*~D+A*B*C*~D+A*B*~C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101111101010111),
    .INIT_LUTF1(16'b1000101010001010),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b1000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2471|picorv32_core/reg0_b12  (
    .a({\picorv32_core/mem_rdata_latched$0$_placeOpt_1 ,_al_u2353_o}),
    .b({_al_u2465_o,_al_u2471_o}),
    .c({\picorv32_core/mem_rdata_latched$1$_placeOpt_3 ,_al_u2470_o}),
    .clk(clk_pad),
    .d({open_n17208,_al_u2468_o}),
    .e({\picorv32_core/mux81_sel_is_1_o ,_al_u2465_o}),
    .f({_al_u2471_o,open_n17224}),
    .q({open_n17228,\picorv32_core/mem_rdata_q [12]}));  // ../src/picorv32.v(508)
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(A*~(0*~B))))"),
    //.LUTF1("(~B*~(D*~(0*~A*~C)))"),
    //.LUTG0("~(~D*~(C*~(A*~(1*~B))))"),
    //.LUTG1("(~B*~(D*~(1*~A*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111101010000),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b1111111101110000),
    .INIT_LUTG1(16'b0000000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2474|picorv32_core/reg0_b13  (
    .a({_al_u2358_o,_al_u2479_o}),
    .b({_al_u2473_o,_al_u2477_o}),
    .c({_al_u2371_o,_al_u1569_o}),
    .clk(clk_pad),
    .d({_al_u1569_o,_al_u2474_o}),
    .e({\picorv32_core/mem_rdata_latched$1$_placeOpt_1 ,_al_u1536_o}),
    .f({_al_u2474_o,open_n17245}),
    .q({open_n17249,\picorv32_core/mem_rdata_q [13]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D)*~(C)*~(B)*A*~(0)+D*~(C)*~(B)*A*~(0)+D*~(C)*B*A*~(0)+D*C*B*A*~(0)+~(D)*~(C)*~(B)*~(A)*0+D*~(C)*~(B)*~(A)*0+~(D)*C*~(B)*~(A)*0+D*C*~(B)*~(A)*0+D*~(C)*B*~(A)*0+D*C*B*~(A)*0+~(D)*~(C)*~(B)*A*0+D*~(C)*~(B)*A*0+~(D)*C*~(B)*A*0+D*C*~(B)*A*0+D*~(C)*B*A*0+D*C*B*A*0)"),
    //.LUT1("(~(D)*~(C)*~(A)*B*~(1)+D*~(C)*~(A)*B*~(1)+D*~(C)*A*B*~(1)+D*C*A*B*~(1)+~(D)*~(C)*~(A)*~(B)*1+D*~(C)*~(A)*~(B)*1+~(D)*C*~(A)*~(B)*1+D*C*~(A)*~(B)*1+D*~(C)*A*~(B)*1+D*C*A*~(B)*1+~(D)*~(C)*~(A)*B*1+D*~(C)*~(A)*B*1+~(D)*C*~(A)*B*1+D*C*~(A)*B*1+D*~(C)*A*B*1+D*C*A*B*1)"),
    .INIT_LUT0(16'b1000101000000010),
    .INIT_LUT1(16'b1111111101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2475 (
    .a({\picorv32_core/mem_rdata_latched [12],_al_u1444_o}),
    .b({_al_u1444_o,\picorv32_core/mem_rdata_latched [12]}),
    .c({\picorv32_core/mem_rdata_latched [6],\picorv32_core/mem_rdata_latched [6]}),
    .d({_al_u2473_o,_al_u2473_o}),
    .mi({open_n17262,_al_u1485_o_placeOpt_2}),
    .fx({open_n17267,_al_u2475_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A*~D)*~(~0*~C*B))"),
    //.LUTF1("0"),
    //.LUTG0("(~(A*~D)*~(~1*~C*B))"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*~C*D+A*B*~C*D"),
    .INIT_LUTF0(16'b1111001101010001),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111111101010101),
    .INIT_LUTG1(16'b0000110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2476|_al_u2477  (
    .a({open_n17270,_al_u2476_o}),
    .b({_al_u1464_o,_al_u2405_o}),
    .c({_al_u1483_o_placeOpt_1,_al_u1579_o}),
    .d({open_n17273,_al_u2475_o}),
    .e({_al_u1481_o_placeOpt_1,_al_u1481_o_placeOpt_1}),
    .f({_al_u2476_o,_al_u2477_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~C*A*D)"),
    //.LUT1("(~(D)*C*~(A)*~(B)+D*C*~(A)*~(B)+~(D)*~(C)*A*~(B)+D*~(C)*A*~(B)+~(D)*C*A*~(B)+D*C*A*~(B)+~(D)*~(C)*~(A)*B+~(D)*C*~(A)*B)"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b0011001001110110),
    .MODE("LOGIC"))
    \_al_u2478|_al_u2292  (
    .a({\picorv32_core/mem_rdata_latched$1$_placeOpt_1 ,\picorv32_core/mem_rdata_latched [2]}),
    .b({\picorv32_core/mem_rdata_latched$0$_placeOpt_1 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_1 }),
    .c({_al_u2291_o,\picorv32_core/mem_rdata_latched$1$_placeOpt_1 }),
    .d({\picorv32_core/mux81_sel_is_1_o ,_al_u2291_o}),
    .f({_al_u2478_o,_al_u2292_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+C*B*~A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("~A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG0("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*~A*D+C*~B*~A*D"),
    //.LUTG1("~A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+~A*B*~D*C+A*B*~D*C+~A*~B*D*C+~A*B*D*C+A*B*D*C"),
    .INIT_LUTF0(16'b1101110111011101),
    .INIT_LUTF1(16'b1101110100000000),
    .INIT_LUTG0(16'b0001000100010001),
    .INIT_LUTG1(16'b1101110111011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2479|_al_u2473  (
    .a({_al_u1597_o,\picorv32_core/mem_rdata_q [13]}),
    .b({\picorv32_core/mem_rdata_latched$0$_placeOpt_1 ,\picorv32_core/mem_xfer_placeOpt_2 }),
    .d({_al_u2473_o,open_n17318}),
    .e({_al_u2478_o,_al_u1485_o_placeOpt_2}),
    .f({_al_u2479_o,_al_u2473_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*D)"),
    //.LUT1("(~A)"),
    .INIT_LUT0(16'b1100110000000000),
    .INIT_LUT1(16'b0101010101010101),
    .MODE("LOGIC"))
    \_al_u2483|_al_u1207  (
    .a({\picorv32_core/latched_compr ,open_n17339}),
    .b({open_n17340,_al_u1206_o}),
    .d({open_n17345,_al_u1204_o}),
    .f({\picorv32_core/n449 [2],_al_u1207_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A)"),
    //.LUT1("(~C)"),
    .INIT_LUT0(16'b0101000001010000),
    .INIT_LUT1(16'b0000111100001111),
    .MODE("LOGIC"))
    \_al_u2484|_al_u1918  (
    .a({open_n17364,_al_u1183_o}),
    .c({mem_la_wdata[0],\picorv32_core/mem_wordsize [0]}),
    .f({n17[0],_al_u1918_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B)"),
    //.LUTF1("(~B)"),
    //.LUTG0("(~B)"),
    //.LUTG1("(~B)"),
    .INIT_LUTF0(16'b0011001100110011),
    .INIT_LUTF1(16'b0011001100110011),
    .INIT_LUTG0(16'b0011001100110011),
    .INIT_LUTG1(16'b0011001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2485|_al_u2486  (
    .b({mem_la_wdata[1],mem_la_wdata[2]}),
    .f({n17[1],n17[2]}));
  EG_PHY_PAD #(
    //.LOCATION("P34"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u539 (
    .ipad(clk),
    .di(clk_pad));  // ../src/top.v(4)
  EG_PHY_PAD #(
    //.LOCATION("P16"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u540 (
    .ipad(resetn_i),
    .di(resetn_i_pad));  // ../src/top.v(5)
  EG_PHY_PAD #(
    //.LOCATION("P13"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u541 (
    .ipad(rxd),
    .di(rxd_pad));  // ../src/top.v(14)
  EG_PHY_PAD #(
    //.LOCATION("P12"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u542 (
    .do({open_n17471,open_n17472,open_n17473,trap_pad}),
    .opad(trap));  // ../src/top.v(6)
  EG_PHY_PAD #(
    //.LOCATION("P14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u543 (
    .do({open_n17488,open_n17489,open_n17490,txd_pad}),
    .opad(txd));  // ../src/top.v(13)
  EG_PHY_MSLICE #(
    //.LUT0("(D*B)"),
    //.LUT1("(D*~C)"),
    .INIT_LUT0(16'b1100110000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u663|_al_u998  (
    .b({open_n17506,\picorv32_core/n663 }),
    .c({\picorv32_core/decoder_pseudo_trigger ,open_n17507}),
    .d({\picorv32_core/decoder_trigger ,\picorv32_core/decoder_trigger }),
    .f({\picorv32_core/n274 ,\picorv32_core/sel39_b0_sel_is_3_o }));
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~B*A*C*~D)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(1*~B*A*C*~D)"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000000000100000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u665|picorv32_core/instr_auipc_reg  (
    .a({open_n17528,\picorv32_core/mem_rdata_latched [4]}),
    .b({open_n17529,\picorv32_core/mem_rdata_latched [3]}),
    .c({open_n17530,_al_u1498_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_auipc ,\picorv32_core/n180 }),
    .e({\picorv32_core/instr_lui ,\picorv32_core/mem_rdata_latched [2]}),
    .f({_al_u665_o,open_n17546}),
    .q({open_n17550,\picorv32_core/instr_auipc }));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~A)"),
    //.LUTF1("(C*A)"),
    //.LUTG0("~(B*~A)"),
    //.LUTG1("(C*A)"),
    .INIT_LUTF0(16'b1011101110111011),
    .INIT_LUTF1(16'b1010000010100000),
    .INIT_LUTG0(16'b1011101110111011),
    .INIT_LUTG1(16'b1010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u669|_al_u753  (
    .a({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .b({open_n17551,resetn_placeOpt_11}),
    .c({\picorv32_core/latched_store ,open_n17552}),
    .f({\picorv32_core/sel15_b0_sel_is_3_o ,\picorv32_core/n447 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~B)"),
    //.LUTF1("(D*B)"),
    //.LUTG0("~(C*~B)"),
    //.LUTG1("(D*B)"),
    .INIT_LUTF0(16'b1100111111001111),
    .INIT_LUTF1(16'b1100110000000000),
    .INIT_LUTG0(16'b1100111111001111),
    .INIT_LUTG1(16'b1100110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u669|_al_u753_placeOpt_1  (
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({open_n17581,resetn_placeOpt_11}),
    .d({\picorv32_core/latched_store ,open_n17584}),
    .f({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,open_n17602}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~B)"),
    //.LUTF1("0"),
    //.LUTG0("~(D*~B)"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1100110011111111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1100110011111111),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u669|_al_u753_placeOpt_2  (
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .d({open_n17614,resetn_placeOpt_11}),
    .e({\picorv32_core/latched_store ,open_n17615}),
    .f({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_2 ,open_n17631}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~B)"),
    //.LUTF1("(D*B)"),
    //.LUTG0("~(A*~B)"),
    //.LUTG1("(D*B)"),
    .INIT_LUTF0(16'b1101110111011101),
    .INIT_LUTF1(16'b1100110000000000),
    .INIT_LUTG0(16'b1101110111011101),
    .INIT_LUTG1(16'b1100110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u669|_al_u753_placeOpt_3  (
    .a({open_n17637,resetn_placeOpt_11}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .d({\picorv32_core/latched_store ,open_n17642}),
    .f({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 ,open_n17660}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~C*B*~D*A+C*B*~D*A+~C*B*D*A+C*B*D*A"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~C*~B*~D*~A+C*~B*~D*~A+~C*B*~D*~A+C*B*~D*~A+~C*~B*D*~A+C*~B*D*~A+~C*B*D*~A+C*B*D*~A+~C*B*~D*A+C*B*~D*A+~C*B*D*A+C*B*D*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1101110111011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u670|picorv32_core/reg17_b9  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({\picorv32_core/reg_out [9],\picorv32_core/latched_stalu }),
    .c({open_n17666,\picorv32_core/reg_out [9]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({open_n17667,\picorv32_core/alu_out_q [9]}),
    .e({\picorv32_core/reg_next_pc [9],\picorv32_core/reg_next_pc [9]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [9],\picorv32_core/n500 [9]}),
    .q({open_n17685,\picorv32_core/reg_pc [9]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*B*~C*~D+~A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*B*~C*~D+~A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1110111001000100),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1110111001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u671|picorv32_core/reg17_b8  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o ,\picorv32_core/sel15_b0_sel_is_3_o }),
    .b({\picorv32_core/reg_next_pc [8],\picorv32_core/latched_stalu }),
    .c({open_n17686,\picorv32_core/reg_out [8]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [8],\picorv32_core/alu_out_q [8]}),
    .e({open_n17687,\picorv32_core/reg_next_pc [8]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [8],\picorv32_core/n500 [8]}),
    .q({open_n17705,\picorv32_core/reg_pc [8]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("A*~B*~D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+A*~B*~D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("A*~B*~D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+A*~B*~D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1110111000100010),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1110111000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u672|picorv32_core/reg17_b7  (
    .a({\picorv32_core/reg_next_pc [7],\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/latched_stalu }),
    .c({open_n17706,\picorv32_core/reg_out [7]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [7],\picorv32_core/alu_out_q [7]}),
    .e({open_n17707,\picorv32_core/reg_next_pc [7]}),
    .sr(resetn),
    .f({\picorv32_core/next_pc [7],\picorv32_core/n500 [7]}),
    .q({open_n17725,\picorv32_core/reg_pc [7]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~D*B*~C*A+D*B*~C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*B*~C*A+D*B*~C*A+~D*B*C*A+D*B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1101110111011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u673|picorv32_core/reg17_b6  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({\picorv32_core/reg_out [6],\picorv32_core/latched_stalu }),
    .c({open_n17726,\picorv32_core/reg_out [6]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({open_n17727,\picorv32_core/alu_out_q [6]}),
    .e({\picorv32_core/reg_next_pc [6],\picorv32_core/reg_next_pc [6]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [6],\picorv32_core/n500 [6]}),
    .q({open_n17745,\picorv32_core/reg_pc [6]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1100110000000000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1100110011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u674|picorv32_core/reg17_b5  (
    .a({open_n17746,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({\picorv32_core/reg_out [5],\picorv32_core/latched_stalu }),
    .c({open_n17747,\picorv32_core/reg_out [5]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/alu_out_q [5]}),
    .e({\picorv32_core/reg_next_pc [5],\picorv32_core/reg_next_pc [5]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [5],\picorv32_core/n500 [5]}),
    .q({open_n17765,\picorv32_core/reg_pc [5]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u675|picorv32_core/reg17_b4  (
    .a({open_n17766,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/latched_stalu }),
    .c({\picorv32_core/reg_next_pc [4],\picorv32_core/reg_out [4]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [4],\picorv32_core/alu_out_q [4]}),
    .e({open_n17767,\picorv32_core/reg_next_pc [4]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [4],\picorv32_core/n500 [4]}),
    .q({open_n17785,\picorv32_core/reg_pc [4]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~B*D*~C*A+B*D*~C*A+~B*D*C*A+B*D*C*A"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~B*~D*~C*~A+B*~D*~C*~A+~B*D*~C*~A+B*D*~C*~A+~B*~D*C*~A+B*~D*C*~A+~B*D*C*~A+B*D*C*~A+~B*D*~C*A+B*D*~C*A+~B*D*C*A+B*D*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1111111101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u676|picorv32_core/reg17_b31  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 }),
    .b({open_n17786,\picorv32_core/latched_stalu }),
    .c({open_n17787,\picorv32_core/reg_out [31]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [31],\picorv32_core/alu_out_q [31]}),
    .e({\picorv32_core/reg_next_pc [31],\picorv32_core/reg_next_pc [31]}),
    .sr(resetn_placeOpt_10),
    .f({\picorv32_core/next_pc [31],\picorv32_core/n500 [31]}),
    .q({open_n17805,\picorv32_core/reg_pc [31]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~C*A*~D*B+C*A*~D*B+~C*A*D*B+C*A*D*B"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~C*~A*~D*~B+C*~A*~D*~B+~C*A*~D*~B+C*A*~D*~B+~C*~A*D*~B+C*~A*D*~B+~C*A*D*~B+C*A*D*~B+~C*A*~D*B+C*A*~D*B+~C*A*D*B+C*A*D*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1011101110111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u677|picorv32_core/reg17_b30  (
    .a({\picorv32_core/reg_out [30],\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 }),
    .b({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 ,\picorv32_core/latched_stalu }),
    .c({open_n17806,\picorv32_core/reg_out [30]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({open_n17807,\picorv32_core/alu_out_q [30]}),
    .e({\picorv32_core/reg_next_pc [30],\picorv32_core/reg_next_pc [30]}),
    .sr(resetn_placeOpt_10),
    .f({\picorv32_core/next_pc [30],\picorv32_core/n500 [30]}),
    .q({open_n17825,\picorv32_core/reg_pc [30]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1100110010101010),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1100110010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u678|picorv32_core/reg17_b3  (
    .a({\picorv32_core/reg_next_pc [3],\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({\picorv32_core/reg_out [3],\picorv32_core/latched_stalu }),
    .c({open_n17826,\picorv32_core/reg_out [3]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/alu_out_q [3]}),
    .e({open_n17827,\picorv32_core/reg_next_pc [3]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [3],\picorv32_core/n500 [3]}),
    .q({open_n17845,\picorv32_core/reg_pc [3]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~C*B*~D*A+C*B*~D*A+~C*B*D*A+C*B*D*A"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~C*~B*~D*~A+C*~B*~D*~A+~C*B*~D*~A+C*B*~D*~A+~C*~B*D*~A+C*~B*D*~A+~C*B*D*~A+C*B*D*~A+~C*B*~D*A+C*B*~D*A+~C*B*D*A+C*B*D*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1101110111011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u679|picorv32_core/reg17_b29  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_2 ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_2 }),
    .b({\picorv32_core/reg_out [29],\picorv32_core/latched_stalu }),
    .c({open_n17846,\picorv32_core/reg_out [29]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({open_n17847,\picorv32_core/alu_out_q [29]}),
    .e({\picorv32_core/reg_next_pc [29],\picorv32_core/reg_next_pc [29]}),
    .sr(resetn_placeOpt_10),
    .f({\picorv32_core/next_pc [29],\picorv32_core/n500 [29]}),
    .q({open_n17865,\picorv32_core/reg_pc [29]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1010101011001100),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1010101011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u680|picorv32_core/reg17_b28  (
    .a({\picorv32_core/reg_out [28],\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 }),
    .b({\picorv32_core/reg_next_pc [28],\picorv32_core/latched_stalu }),
    .c({open_n17866,\picorv32_core/reg_out [28]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 ,\picorv32_core/alu_out_q [28]}),
    .e({open_n17867,\picorv32_core/reg_next_pc [28]}),
    .sr(resetn_placeOpt_10),
    .f({\picorv32_core/next_pc [28],\picorv32_core/n500 [28]}),
    .q({open_n17885,\picorv32_core/reg_pc [28]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~D*B*~C*A+D*B*~C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*B*~C*A+D*B*~C*A+~D*B*C*A+D*B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1101110111011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u681|picorv32_core/reg17_b27  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_2 ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_2 }),
    .b({\picorv32_core/reg_out [27],\picorv32_core/latched_stalu }),
    .c({open_n17886,\picorv32_core/reg_out [27]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({open_n17887,\picorv32_core/alu_out_q [27]}),
    .e({\picorv32_core/reg_next_pc [27],\picorv32_core/reg_next_pc [27]}),
    .sr(resetn),
    .f({\picorv32_core/next_pc [27],\picorv32_core/n500 [27]}),
    .q({open_n17905,\picorv32_core/reg_pc [27]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~C*A*~D*B+C*A*~D*B+~C*A*D*B+C*A*D*B"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~C*~A*~D*~B+C*~A*~D*~B+~C*A*~D*~B+C*A*~D*~B+~C*~A*D*~B+C*~A*D*~B+~C*A*D*~B+C*A*D*~B+~C*A*~D*B+C*A*~D*B+~C*A*D*B+C*A*D*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1011101110111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u682|picorv32_core/reg17_b26  (
    .a({\picorv32_core/reg_out [26],\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_2 }),
    .b({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_2 ,\picorv32_core/latched_stalu }),
    .c({open_n17906,\picorv32_core/reg_out [26]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({open_n17907,\picorv32_core/alu_out_q [26]}),
    .e({\picorv32_core/reg_next_pc [26],\picorv32_core/reg_next_pc [26]}),
    .sr(resetn),
    .f({\picorv32_core/next_pc [26],\picorv32_core/n500 [26]}),
    .q({open_n17925,\picorv32_core/reg_pc [26]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u683|picorv32_core/reg17_b25  (
    .a({open_n17926,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 }),
    .b({\picorv32_core/reg_next_pc [25],\picorv32_core/latched_stalu }),
    .c({\picorv32_core/reg_out [25],\picorv32_core/reg_out [25]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 ,\picorv32_core/alu_out_q [25]}),
    .e({open_n17927,\picorv32_core/reg_next_pc [25]}),
    .sr(resetn_placeOpt_10),
    .f({\picorv32_core/next_pc [25],\picorv32_core/n500 [25]}),
    .q({open_n17945,\picorv32_core/reg_pc [25]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("A*~B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("A*~B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1110001011100010),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1110001011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u684|picorv32_core/reg17_b24  (
    .a({\picorv32_core/reg_next_pc [24],\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 }),
    .b({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 ,\picorv32_core/latched_stalu }),
    .c({\picorv32_core/reg_out [24],\picorv32_core/reg_out [24]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({open_n17946,\picorv32_core/alu_out_q [24]}),
    .e({open_n17947,\picorv32_core/reg_next_pc [24]}),
    .sr(resetn_placeOpt_10),
    .f({\picorv32_core/next_pc [24],\picorv32_core/n500 [24]}),
    .q({open_n17965,\picorv32_core/reg_pc [24]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~C*D*~B*A+C*D*~B*A+~C*D*B*A+C*D*B*A"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~C*~D*~B*~A+C*~D*~B*~A+~C*D*~B*~A+C*D*~B*~A+~C*~D*B*~A+C*~D*B*~A+~C*D*B*~A+C*D*B*~A+~C*D*~B*A+C*D*~B*A+~C*D*B*A+C*D*B*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1111111101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u685|picorv32_core/reg17_b23  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_2 ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_2 }),
    .b({open_n17966,\picorv32_core/latched_stalu }),
    .c({open_n17967,\picorv32_core/reg_out [23]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [23],\picorv32_core/alu_out_q [23]}),
    .e({\picorv32_core/reg_next_pc [23],\picorv32_core/reg_next_pc [23]}),
    .sr(resetn),
    .f({\picorv32_core/next_pc [23],\picorv32_core/n500 [23]}),
    .q({open_n17985,\picorv32_core/reg_pc [23]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*B*~D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*B*~D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*B*~D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*B*~D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1110111001000100),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1110111001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u686|picorv32_core/reg17_b22  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 }),
    .b({\picorv32_core/reg_next_pc [22],\picorv32_core/latched_stalu }),
    .c({open_n17986,\picorv32_core/reg_out [22]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [22],\picorv32_core/alu_out_q [22]}),
    .e({open_n17987,\picorv32_core/reg_next_pc [22]}),
    .sr(resetn_placeOpt_10),
    .f({\picorv32_core/next_pc [22],\picorv32_core/n500 [22]}),
    .q({open_n18005,\picorv32_core/reg_pc [22]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b0101010100000000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1111111110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u687|picorv32_core/reg17_b21  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 }),
    .b({open_n18006,\picorv32_core/latched_stalu }),
    .c({open_n18007,\picorv32_core/reg_out [21]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/reg_next_pc [21],\picorv32_core/alu_out_q [21]}),
    .e({\picorv32_core/reg_out [21],\picorv32_core/reg_next_pc [21]}),
    .sr(resetn_placeOpt_10),
    .f({\picorv32_core/next_pc [21],\picorv32_core/n500 [21]}),
    .q({open_n18025,\picorv32_core/reg_pc [21]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*B*~C*~D+~A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*B*~C*~D+~A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1110111001000100),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1110111001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u688|picorv32_core/reg17_b20  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o ,\picorv32_core/sel15_b0_sel_is_3_o }),
    .b({\picorv32_core/reg_next_pc [20],\picorv32_core/latched_stalu }),
    .c({open_n18026,\picorv32_core/reg_out [20]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [20],\picorv32_core/alu_out_q [20]}),
    .e({open_n18027,\picorv32_core/reg_next_pc [20]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [20],\picorv32_core/n500 [20]}),
    .q({open_n18045,\picorv32_core/reg_pc [20]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("A*~B*~C*~D+A*~B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("A*~B*~C*~D+A*~B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1110111000100010),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1110111000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u689|picorv32_core/reg17_b2  (
    .a({\picorv32_core/reg_next_pc [2],\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/latched_stalu }),
    .c({open_n18046,\picorv32_core/reg_out [2]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [2],\picorv32_core/alu_out_q [2]}),
    .e({open_n18047,\picorv32_core/reg_next_pc [2]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [2],\picorv32_core/n500 [2]}),
    .q({open_n18065,\picorv32_core/reg_pc [2]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1111010110100000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1111010110100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u690|picorv32_core/reg17_b19  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_3 }),
    .b({open_n18066,\picorv32_core/latched_stalu }),
    .c({\picorv32_core/reg_out [19],\picorv32_core/reg_out [19]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/reg_next_pc [19],\picorv32_core/alu_out_q [19]}),
    .e({open_n18067,\picorv32_core/reg_next_pc [19]}),
    .sr(resetn_placeOpt_10),
    .f({\picorv32_core/next_pc [19],\picorv32_core/n500 [19]}),
    .q({open_n18085,\picorv32_core/reg_pc [19]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*C*~B*~D+A*C*~B*~D+~A*C*B*~D+A*C*B*~D+A*~C*~B*D+A*C*~B*D+A*~C*B*D+A*C*B*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*C*~B*~D+A*C*~B*~D+~A*C*B*~D+A*C*B*~D+A*~C*~B*D+A*C*~B*D+A*~C*B*D+A*C*B*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1010101011110000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1010101011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u691|picorv32_core/reg17_b18  (
    .a({\picorv32_core/reg_out [18],\picorv32_core/sel15_b0_sel_is_3_o }),
    .b({open_n18086,\picorv32_core/latched_stalu }),
    .c({\picorv32_core/reg_next_pc [18],\picorv32_core/reg_out [18]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/sel15_b0_sel_is_3_o ,\picorv32_core/alu_out_q [18]}),
    .e({open_n18087,\picorv32_core/reg_next_pc [18]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [18],\picorv32_core/n500 [18]}),
    .q({open_n18105,\picorv32_core/reg_pc [18]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*~B*C*~D+~A*B*C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*~B*C*~D+~A*B*C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1111101001010000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1111101001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u692|picorv32_core/reg17_b17  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({open_n18106,\picorv32_core/latched_stalu }),
    .c({\picorv32_core/reg_next_pc [17],\picorv32_core/reg_out [17]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [17],\picorv32_core/alu_out_q [17]}),
    .e({open_n18107,\picorv32_core/reg_next_pc [17]}),
    .sr(resetn),
    .f({\picorv32_core/next_pc [17],\picorv32_core/n500 [17]}),
    .q({open_n18125,\picorv32_core/reg_pc [17]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1111000010101010),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1111000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u693|picorv32_core/reg17_b16  (
    .a({\picorv32_core/reg_next_pc [16],\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({open_n18126,\picorv32_core/latched_stalu }),
    .c({\picorv32_core/reg_out [16],\picorv32_core/reg_out [16]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/alu_out_q [16]}),
    .e({open_n18127,\picorv32_core/reg_next_pc [16]}),
    .sr(resetn),
    .f({\picorv32_core/next_pc [16],\picorv32_core/n500 [16]}),
    .q({open_n18145,\picorv32_core/reg_pc [16]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~C*A*~B*D+C*A*~B*D+~C*A*B*D+C*A*B*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~C*~A*~B*~D+C*~A*~B*~D+~C*A*~B*~D+C*A*~B*~D+~C*~A*B*~D+C*~A*B*~D+~C*A*B*~D+C*A*B*~D+~C*A*~B*D+C*A*~B*D+~C*A*B*D+C*A*B*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1010101011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u694|picorv32_core/reg17_b15  (
    .a({\picorv32_core/reg_out [15],\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({open_n18146,\picorv32_core/latched_stalu }),
    .c({open_n18147,\picorv32_core/reg_out [15]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/alu_out_q [15]}),
    .e({\picorv32_core/reg_next_pc [15],\picorv32_core/reg_next_pc [15]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [15],\picorv32_core/n500 [15]}),
    .q({open_n18165,\picorv32_core/reg_pc [15]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~D*B*~C*A+D*B*~C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*B*~C*A+D*B*~C*A+~D*B*C*A+D*B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1101110111011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u695|picorv32_core/reg17_b14  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({\picorv32_core/reg_out [14],\picorv32_core/latched_stalu }),
    .c({open_n18166,\picorv32_core/reg_out [14]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({open_n18167,\picorv32_core/alu_out_q [14]}),
    .e({\picorv32_core/reg_next_pc [14],\picorv32_core/reg_next_pc [14]}),
    .sr(resetn),
    .f({\picorv32_core/next_pc [14],\picorv32_core/n500 [14]}),
    .q({open_n18185,\picorv32_core/reg_pc [14]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u696|picorv32_core/reg17_b13  (
    .a({open_n18186,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({\picorv32_core/reg_out [13],\picorv32_core/latched_stalu }),
    .c({\picorv32_core/reg_next_pc [13],\picorv32_core/reg_out [13]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/alu_out_q [13]}),
    .e({open_n18187,\picorv32_core/reg_next_pc [13]}),
    .sr(resetn),
    .f({\picorv32_core/next_pc [13],\picorv32_core/n500 [13]}),
    .q({open_n18205,\picorv32_core/reg_pc [13]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1010101011110000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1010101011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u697|picorv32_core/reg17_b12  (
    .a({\picorv32_core/reg_out [12],\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({open_n18206,\picorv32_core/latched_stalu }),
    .c({\picorv32_core/reg_next_pc [12],\picorv32_core/reg_out [12]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/alu_out_q [12]}),
    .e({open_n18207,\picorv32_core/reg_next_pc [12]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [12],\picorv32_core/n500 [12]}),
    .q({open_n18225,\picorv32_core/reg_pc [12]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~A*~B*C*~D+~A*B*C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~A*~B*C*~D+~A*B*C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1111101001010000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1111101001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u698|picorv32_core/reg17_b11  (
    .a({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({open_n18226,\picorv32_core/latched_stalu }),
    .c({\picorv32_core/reg_next_pc [11],\picorv32_core/reg_out [11]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/reg_out [11],\picorv32_core/alu_out_q [11]}),
    .e({open_n18227,\picorv32_core/reg_next_pc [11]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [11],\picorv32_core/n500 [11]}),
    .q({open_n18245,\picorv32_core/reg_pc [11]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(0)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+0*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTF1("~C*A*~D*B+C*A*~D*B+~C*A*D*B+C*A*D*B"),
    //.LUTG0("(1*~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*~(A)+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)+~(1)*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A+1*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A)"),
    //.LUTG1("~C*~A*~D*~B+C*~A*~D*~B+~C*A*~D*~B+C*A*~D*~B+~C*~A*D*~B+C*~A*D*~B+~C*A*D*~B+C*A*D*~B+~C*A*~D*B+C*A*~D*B+~C*A*D*B+C*A*D*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1111110101110101),
    .INIT_LUTG1(16'b1011101110111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u699|picorv32_core/reg17_b10  (
    .a({\picorv32_core/reg_out [10],\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 }),
    .b({\picorv32_core/sel15_b0_sel_is_3_o_placeOpt_1 ,\picorv32_core/latched_stalu }),
    .c({open_n18246,\picorv32_core/reg_out [10]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({open_n18247,\picorv32_core/alu_out_q [10]}),
    .e({\picorv32_core/reg_next_pc [10],\picorv32_core/reg_next_pc [10]}),
    .sr(resetn_placeOpt_7),
    .f({\picorv32_core/next_pc [10],\picorv32_core/n500 [10]}),
    .q({open_n18265,\picorv32_core/reg_pc [10]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D"),
    //.LUTG0("(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1110111000100010),
    .INIT_LUTF1(16'b0000000010101010),
    .INIT_LUTG0(16'b1110111000100010),
    .INIT_LUTG1(16'b1111111110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u701|_al_u710  (
    .a({\picorv32_core/n30 [7],\picorv32_core/n30 [8]}),
    .b({open_n18266,_al_u700_o}),
    .d({_al_u700_o,\picorv32_core/pcpi_rs1$10$ }),
    .e({\picorv32_core/pcpi_rs1$9$ ,open_n18271}),
    .f({mem_la_addr[9],mem_la_addr[10]}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b1010111110100000),
    .MODE("LOGIC"))
    \_al_u703|_al_u706  (
    .a({\picorv32_core/pcpi_rs1$7$ ,open_n18292}),
    .b({open_n18293,\picorv32_core/pcpi_rs1$4$ }),
    .c({_al_u700_o,_al_u700_o}),
    .d({\picorv32_core/n30 [5],\picorv32_core/n30 [2]}),
    .f({mem_la_addr[7],mem_la_addr[4]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~C*~D)*~((~0*~A))*~(B)+(~C*~D)*(~0*~A)*~(B)+~((~C*~D))*(~0*~A)*B+(~C*~D)*(~0*~A)*B)"),
    //.LUTF1("A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("~((~C*~D)*~((~1*~A))*~(B)+(~C*~D)*(~1*~A)*~(B)+~((~C*~D))*(~1*~A)*B+(~C*~D)*(~1*~A)*B)"),
    //.LUTG1("A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1011101110111000),
    .INIT_LUTF1(16'b1010111110100000),
    .INIT_LUTG0(16'b1111111111111100),
    .INIT_LUTG1(16'b1010111110100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u705|_al_u1171  (
    .a({\picorv32_core/pcpi_rs1$5$ ,\picorv32_core/pcpi_rs1$5$ }),
    .b({open_n18314,_al_u700_o}),
    .c({_al_u700_o,\picorv32_core/n30 [3]}),
    .d({\picorv32_core/n30 [3],\picorv32_core/n30 [4]}),
    .e({open_n18317,\picorv32_core/pcpi_rs1$6$ }),
    .f({mem_la_addr[5],\eq2/or_xor_i0$1$_i1$1$_o_o_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    //.LUTF1("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    //.LUTG0("(1*C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    //.LUTG1("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1110111001000100),
    .INIT_LUTG0(16'b1101000010000000),
    .INIT_LUTG1(16'b1110111001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u707|_al_u816  (
    .a({_al_u700_o_placeOpt_1,_al_u700_o_placeOpt_1}),
    .b({\picorv32_core/n30 [1],\picorv32_core/pcpi_rs1$3$ }),
    .c({open_n18338,mem_la_addr[2]}),
    .d({\picorv32_core/pcpi_rs1$3$ ,\picorv32_core/n30 [1]}),
    .e({open_n18341,\uart/uart_status_rx }),
    .f({mem_la_addr[3],_al_u816_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~C*D)*~((0*~A))*~(B)+(~C*D)*(0*~A)*~(B)+~((~C*D))*(0*~A)*B+(~C*D)*(0*~A)*B)"),
    //.LUTF1("D*~B*~A*~C+D*~B*A*~C+D*~B*~A*C+D*~B*A*C"),
    //.LUTG0("~((~C*D)*~((1*~A))*~(B)+(~C*D)*(1*~A)*~(B)+~((~C*D))*(1*~A)*B+(~C*D)*(1*~A)*B)"),
    //.LUTG1("D*~B*~A*~C+~D*B*~A*~C+D*B*~A*~C+D*~B*A*~C+~D*B*A*~C+D*B*A*~C+D*~B*~A*C+~D*B*~A*C+D*B*~A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b0011001100000000),
    .INIT_LUTG0(16'b1011100010111011),
    .INIT_LUTG1(16'b1111111111001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u708|_al_u812  (
    .a({open_n18362,\picorv32_core/pcpi_rs1$2$ }),
    .b({_al_u700_o_placeOpt_1,_al_u700_o_placeOpt_1}),
    .c({open_n18363,\picorv32_core/n30 [0]}),
    .d({\picorv32_core/n30 [0],\picorv32_core/n30 [1]}),
    .e({\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$3$ }),
    .f({mem_la_addr[2],_al_u812_o}));
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0101111101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg  (
    .a({initial_reset[1],open_n18386}),
    .c({initial_reset[0],resetn_i_pad}),
    .clk(clk_pad),
    .d({open_n18390,\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .f({\eq0/or_xor_i0$0$_i1$0$_o_o ,open_n18404}),
    .q({open_n18408,resetn}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~B)"),
    //.LUT1("~(A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001000100010),
    .INIT_LUT1(16'b0101010111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_1  (
    .a({initial_reset[1],resetn_i_pad}),
    .b({open_n18409,\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .clk(clk_pad),
    .d({initial_reset[0],open_n18413}),
    .q({open_n18432,resetn_placeOpt_1}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0011001111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_10  (
    .b({initial_reset[1],open_n18435}),
    .c({open_n18436,resetn_i_pad}),
    .clk(clk_pad),
    .d({initial_reset[0],\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .q({open_n18456,resetn_placeOpt_10}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A)"),
    //.LUT1("~(D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010001000100),
    .INIT_LUT1(16'b0000111111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_11  (
    .a({open_n18457,\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .b({open_n18458,resetn_i_pad}),
    .c({initial_reset[0],open_n18459}),
    .clk(clk_pad),
    .d({initial_reset[1],open_n18461}),
    .q({open_n18480,resetn_placeOpt_11}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~B)"),
    //.LUT1("~(A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001000100010),
    .INIT_LUT1(16'b0101010111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_12  (
    .a({initial_reset[1],resetn_i_pad}),
    .b({open_n18481,\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .clk(clk_pad),
    .d({initial_reset[0],open_n18485}),
    .q({open_n18504,resetn_placeOpt_12}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A)"),
    //.LUT1("~(B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000001010000),
    .INIT_LUT1(16'b0111011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_13  (
    .a({initial_reset[0],\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .b({initial_reset[1],open_n18505}),
    .c({open_n18506,resetn_i_pad}),
    .clk(clk_pad),
    .q({open_n18528,resetn_placeOpt_13}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A)"),
    //.LUT1("~(C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010001000100),
    .INIT_LUT1(16'b0011111100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_14  (
    .a({open_n18529,\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .b({initial_reset[0],resetn_i_pad}),
    .c({initial_reset[1],open_n18530}),
    .clk(clk_pad),
    .q({open_n18552,resetn_placeOpt_14}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A)"),
    //.LUT1("~(B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010001000100),
    .INIT_LUT1(16'b0011001111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_15  (
    .a({open_n18553,\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .b({initial_reset[1],resetn_i_pad}),
    .clk(clk_pad),
    .d({initial_reset[0],open_n18557}),
    .q({open_n18576,resetn_placeOpt_15}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~B)"),
    //.LUT1("~(A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001100000000),
    .INIT_LUT1(16'b0101010111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_16  (
    .a({initial_reset[1],open_n18577}),
    .b({open_n18578,\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .clk(clk_pad),
    .d({initial_reset[0],resetn_i_pad}),
    .q({open_n18600,resetn_placeOpt_16}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A)"),
    //.LUT1("~(A*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010001000100),
    .INIT_LUT1(16'b0111011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_17  (
    .a({initial_reset[1],\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .b({initial_reset[0],resetn_i_pad}),
    .clk(clk_pad),
    .q({open_n18624,resetn_placeOpt_17}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A)"),
    //.LUT1("~(A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010001000100),
    .INIT_LUT1(16'b0101010111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_2  (
    .a({initial_reset[1],\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .b({open_n18625,resetn_i_pad}),
    .clk(clk_pad),
    .d({initial_reset[0],open_n18629}),
    .q({open_n18648,resetn_placeOpt_2}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A)"),
    //.LUT1("~(B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000001010000),
    .INIT_LUT1(16'b0011001111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_3  (
    .a({open_n18649,\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .b({initial_reset[1],open_n18650}),
    .c({open_n18651,resetn_i_pad}),
    .clk(clk_pad),
    .d({initial_reset[0],open_n18653}),
    .q({open_n18672,resetn_placeOpt_3}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~D)"),
    //.LUT1("~(B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b0011111100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_4  (
    .a({open_n18673,resetn_i_pad}),
    .b({initial_reset[1],open_n18674}),
    .c({initial_reset[0],open_n18675}),
    .clk(clk_pad),
    .d({open_n18677,\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .q({open_n18696,resetn_placeOpt_4}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A)"),
    //.LUT1("~(B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010001000100),
    .INIT_LUT1(16'b0011001111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_5  (
    .a({open_n18697,\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .b({initial_reset[1],resetn_i_pad}),
    .clk(clk_pad),
    .d({initial_reset[0],open_n18701}),
    .q({open_n18720,resetn_placeOpt_5}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A)"),
    //.LUT1("~(A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010001000100),
    .INIT_LUT1(16'b0101010111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_6  (
    .a({initial_reset[1],\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .b({open_n18721,resetn_i_pad}),
    .clk(clk_pad),
    .d({initial_reset[0],open_n18725}),
    .q({open_n18744,resetn_placeOpt_6}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~D)"),
    //.LUT1("~(A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001100),
    .INIT_LUT1(16'b0101010111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_7  (
    .a({initial_reset[1],open_n18745}),
    .b({open_n18746,resetn_i_pad}),
    .clk(clk_pad),
    .d({initial_reset[0],\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .q({open_n18768,resetn_placeOpt_7}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~D)"),
    //.LUT1("~(C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001100),
    .INIT_LUT1(16'b0011111100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_8  (
    .b({initial_reset[0],resetn_i_pad}),
    .c({initial_reset[1],open_n18771}),
    .clk(clk_pad),
    .d({open_n18773,\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .q({open_n18792,resetn_placeOpt_8}));  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~A)"),
    //.LUT1("~(D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010100000000),
    .INIT_LUT1(16'b0011001111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u752|resetn_reg_placeOpt_9  (
    .a({open_n18793,\eq0/or_xor_i0$0$_i1$0$_o_o }),
    .b({initial_reset[0],open_n18794}),
    .clk(clk_pad),
    .d({initial_reset[1],resetn_i_pad}),
    .q({open_n18816,resetn_placeOpt_9}));  // ../src/top.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~D))"),
    //.LUT1("~(C*~B)"),
    .INIT_LUT0(16'b1111000000110000),
    .INIT_LUT1(16'b1100111111001111),
    .MODE("LOGIC"))
    \_al_u754|_al_u1615  (
    .b({trap_pad,trap_pad}),
    .c({resetn_placeOpt_13,resetn_placeOpt_13}),
    .d({open_n18821,\picorv32_core/mem_state [1]}),
    .f({\picorv32_core/n111 ,_al_u1615_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*~C*D+B*~A*~C*D+~B*~A*C*D+B*~A*C*D"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*~A*~C*D+B*~A*~C*D+~B*~A*C*D+B*~A*C*D"),
    //.LUTG0("0"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0101010100000000),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u799|_al_u800  (
    .a(\uart/uart_status_txd [1:0]),
    .d({open_n18846,_al_u799_o}),
    .e({\uart/uart_status_txd [2],\uart/uart_status_txd [3]}),
    .f({_al_u799_o,\uart/n9_lutinv }));
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(B*C*A*D)"),
    //.LUT1("~(~D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u801|uart/uart_trigger_tx_reg  (
    .a({open_n18867,_al_u1168_o}),
    .b({\uart/n9_lutinv ,\uart/n9_lutinv }),
    .c({open_n18868,_al_u1175_o}),
    .ce(\picorv32_core/n524$4$_en_al_n602 ),
    .clk(clk_pad),
    .d({\uart/uart_trigger_tx ,_al_u1179_o}),
    .sr(resetn),
    .f({\uart/n30 ,open_n18881}),
    .q({open_n18885,\uart/uart_trigger_tx }));  // ../src/uart.v(102)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u802|picorv32_core/instr_rdcycle_reg  (
    .b({resetn_placeOpt_8,open_n18888}),
    .c({open_n18889,_al_u1143_o}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/n274 ,_al_u1100_o}),
    .f({\picorv32_core/u449_sel_is_0_o ,open_n18907}),
    .q({open_n18911,\picorv32_core/instr_rdcycle }));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000001100000011),
    .INIT_LUTG0(16'b0000000010101010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u803|_al_u1549  (
    .a({open_n18912,\picorv32_core/n664_lutinv_placeOpt_6 }),
    .b({\picorv32_core/is_alu_reg_imm ,open_n18913}),
    .c({\picorv32_core/is_lb_lh_lw_lbu_lhu ,open_n18914}),
    .d({open_n18917,\picorv32_core/n524 [7]}),
    .e({\picorv32_core/instr_jalr ,\picorv32_core/is_lb_lh_lw_lbu_lhu }),
    .f({_al_u803_o,\picorv32_core/sel40_b0/or_or_B4_B5_o_or_B6__o_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)*~(~0*~C))"),
    //.LUTF1("(~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)*~(~0*~C))"),
    //.LUTG0("(~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)*~(~1*~C))"),
    //.LUTG1("(~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)*~(~1*~C))"),
    .INIT_LUTF0(16'b0010000001110000),
    .INIT_LUTF1(16'b0010000001110000),
    .INIT_LUTG0(16'b0010001001110111),
    .INIT_LUTG1(16'b0010001001110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u810|_al_u815  (
    .a({_al_u700_o,_al_u700_o}),
    .b({\picorv32_core/pcpi_rs1$3$ ,\picorv32_core/pcpi_rs1$3$ }),
    .c({mem_la_addr[2],mem_la_addr[2]}),
    .d({\picorv32_core/n30 [1],\picorv32_core/n30 [1]}),
    .e(\uart/uart_odr [2:1]),
    .f({_al_u810_o,_al_u815_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(0*C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    //.LUT1("(1*C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1101000010000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u811 (
    .a({_al_u700_o_placeOpt_1,_al_u700_o_placeOpt_1}),
    .b({\picorv32_core/pcpi_rs1$3$ ,\picorv32_core/pcpi_rs1$3$ }),
    .c({mem_la_addr[2],mem_la_addr[2]}),
    .d({\picorv32_core/n30 [1],\picorv32_core/n30 [1]}),
    .mi({open_n18972,\uart/uart_status_fe }),
    .fx({open_n18977,_al_u811_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*B*D*~A+~C*B*D*A"),
    //.LUTF1("~C*B*A*~D+C*B*A*~D"),
    //.LUTG0("~C*~B*~D*~A+~C*~B*D*~A+~C*B*D*~A+~C*~B*~D*A+~C*~B*D*A+~C*B*D*A"),
    //.LUTG1("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000000010001000),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b0000000010111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u813|_al_u817  (
    .a({\picorv32_core/pcpi_rs1$2$ ,open_n18980}),
    .b({_al_u700_o_placeOpt_1,_al_u700_o_placeOpt_1}),
    .c({open_n18981,\uart/uart_idr [1]}),
    .d({\uart/uart_idr [2],\picorv32_core/pcpi_rs1$2$ }),
    .e({\picorv32_core/n30 [0],\picorv32_core/n30 [0]}),
    .f({_al_u813_o,_al_u817_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b0000000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u826|picorv32_core/instr_xori_reg  (
    .a({open_n19004,\picorv32_core/is_alu_reg_imm }),
    .b({\picorv32_core/instr_xori ,\picorv32_core/mem_rdata_q [12]}),
    .c({open_n19005,\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_xor ,\picorv32_core/mem_rdata_q [14]}),
    .sr(resetn_placeOpt_8),
    .f({_al_u826_o,open_n19018}),
    .q({open_n19022,\picorv32_core/instr_xori }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(~D*~C)"),
    //.LUTG0("~C*~B*D*A+C*~B*D*A"),
    //.LUTG1("(~D*~C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0010001000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u827|picorv32_core/instr_ori_reg  (
    .a({open_n19023,\picorv32_core/mem_rdata_q [14]}),
    .b({open_n19024,\picorv32_core/mem_rdata_q [12]}),
    .c({\picorv32_core/instr_or ,open_n19025}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_ori ,\picorv32_core/mem_rdata_q [13]}),
    .e({open_n19026,\picorv32_core/is_alu_reg_imm }),
    .sr(resetn_placeOpt_8),
    .f({_al_u827_o,open_n19041}),
    .q({open_n19045,\picorv32_core/instr_ori }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(~D*~A)"),
    //.LUTG0("A*~C*B*D+A*C*B*D"),
    //.LUTG1("(~D*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b1000100000000000),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u828|picorv32_core/instr_andi_reg  (
    .a({\picorv32_core/instr_and ,\picorv32_core/is_alu_reg_imm }),
    .b({open_n19046,\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_andi ,\picorv32_core/mem_rdata_q [14]}),
    .e({open_n19049,\picorv32_core/mem_rdata_q [12]}),
    .sr(resetn_placeOpt_8),
    .f({_al_u828_o,open_n19064}),
    .q({open_n19068,\picorv32_core/instr_andi }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+A*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*B*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*B*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+A*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1)"),
    .INIT_LUT0(16'b0111011100000000),
    .INIT_LUT1(16'b0011011111110111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u833 (
    .a({_al_u826_o,_al_u826_o}),
    .b({_al_u827_o,_al_u827_o}),
    .c({\picorv32_core/pcpi_rs1$11$ ,_al_u828_o}),
    .d({_al_u828_o,\picorv32_core/pcpi_rs1$11$ }),
    .mi({open_n19081,\picorv32_core/pcpi_rs2$11$ }),
    .fx({open_n19086,_al_u833_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(0*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)))"),
    //.LUTF1("~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+~D*~B*C*A+D*~B*C*A+~D*B*C*A"),
    //.LUTG0("~(~D*~(1*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)))"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+~D*~B*C*A+D*~B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b1111111111001010),
    .INIT_LUTG1(16'b0111001101111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u835|picorv32_core/reg14_b12  (
    .a({_al_u828_o,\picorv32_core/n434 [12]}),
    .b({_al_u827_o,\picorv32_core/n433 [12]}),
    .c({\picorv32_core/pcpi_rs2$12$ ,\picorv32_core/instr_sub }),
    .clk(clk_pad),
    .d({_al_u826_o,_al_u835_o}),
    .e({\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u835_o,open_n19105}),
    .q({open_n19109,\picorv32_core/alu_out_q [12]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(0*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)))"),
    //.LUTF1("~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+~D*~B*C*A+D*~B*C*A+~D*B*C*A"),
    //.LUTG0("~(~D*~(1*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)))"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+~D*~B*C*A+D*~B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b1111111111001010),
    .INIT_LUTG1(16'b0111001101111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u837|picorv32_core/reg14_b13  (
    .a({_al_u828_o,\picorv32_core/n434 [13]}),
    .b({_al_u827_o,\picorv32_core/n433 [13]}),
    .c({\picorv32_core/pcpi_rs2$13$ ,\picorv32_core/instr_sub }),
    .clk(clk_pad),
    .d({_al_u826_o,_al_u837_o}),
    .e({\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u837_o,open_n19126}),
    .q({open_n19130,\picorv32_core/alu_out_q [13]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(0*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)))"),
    //.LUTF1("~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D"),
    //.LUTG0("~(~A*~(1*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)))"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b0101111100000000),
    .INIT_LUTG0(16'b1110111011111010),
    .INIT_LUTG1(16'b0011111101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u843|picorv32_core/reg14_b16  (
    .a({_al_u826_o,_al_u843_o}),
    .b({_al_u828_o,\picorv32_core/n433 [16]}),
    .c({_al_u827_o,\picorv32_core/n434 [16]}),
    .clk(clk_pad),
    .d({\picorv32_core/pcpi_rs2$16$ ,\picorv32_core/instr_sub }),
    .e({\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u843_o,open_n19147}),
    .q({open_n19151,\picorv32_core/alu_out_q [16]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(0*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)))"),
    //.LUTF1("(~(D)*~(B)*~(A)*C*~(0)+D*~(B)*~(A)*C*~(0)+~(D)*B*~(A)*C*~(0)+~(D)*~(B)*A*C*~(0)+D*~(B)*A*C*~(0)+~(D)*B*A*C*~(0)+~(D)*~(B)*~(A)*~(C)*0+D*~(B)*~(A)*~(C)*0+~(D)*B*~(A)*~(C)*0+~(D)*~(B)*A*~(C)*0+D*~(B)*A*~(C)*0+~(D)*B*A*~(C)*0+~(D)*~(B)*~(A)*C*0+D*~(B)*~(A)*C*0+~(D)*B*~(A)*C*0+D*B*~(A)*C*0+~(D)*~(B)*A*C*0+D*~(B)*A*C*0)"),
    //.LUTG0("~(~D*~(1*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)))"),
    //.LUTG1("(~(D)*~(B)*~(A)*C*~(1)+D*~(B)*~(A)*C*~(1)+~(D)*B*~(A)*C*~(1)+~(D)*~(B)*A*C*~(1)+D*~(B)*A*C*~(1)+~(D)*B*A*C*~(1)+~(D)*~(B)*~(A)*~(C)*1+D*~(B)*~(A)*~(C)*1+~(D)*B*~(A)*~(C)*1+~(D)*~(B)*A*~(C)*1+D*~(B)*A*~(C)*1+~(D)*B*A*~(C)*1+~(D)*~(B)*~(A)*C*1+D*~(B)*~(A)*C*1+~(D)*B*~(A)*C*1+D*B*~(A)*C*1+~(D)*~(B)*A*C*1+D*~(B)*A*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b1111111111001010),
    .INIT_LUTG1(16'b0111001101111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u845|picorv32_core/reg14_b17  (
    .a({_al_u828_o,\picorv32_core/n434 [17]}),
    .b({_al_u827_o,\picorv32_core/n433 [17]}),
    .c({\picorv32_core/pcpi_rs1$17$ ,\picorv32_core/instr_sub }),
    .clk(clk_pad),
    .d({_al_u826_o,_al_u845_o}),
    .e({\picorv32_core/pcpi_rs2$17$ ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u845_o,open_n19168}),
    .q({open_n19172,\picorv32_core/alu_out_q [17]}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("~D*~C*~B*A+D*~C*~B*A+~D*C*~B*A+~D*~C*B*A+D*~C*B*A+~D*C*B*A"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("~D*~C*~B*~A+D*~C*~B*~A+~D*C*~B*~A+~D*~C*B*~A+D*~C*B*~A+~D*C*B*~A+~D*~C*~B*A+D*~C*~B*A+~D*C*~B*A+D*C*~B*A+~D*~C*B*A+D*~C*B*A"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b0010111101111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u847|_al_u865  (
    .a({\picorv32_core/pcpi_rs2$18$ ,_al_u826_o}),
    .b({_al_u828_o,_al_u827_o}),
    .c({_al_u827_o,_al_u828_o}),
    .d({_al_u826_o,\picorv32_core/pcpi_rs1$26$ }),
    .e({\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs2$26$ }),
    .f({_al_u847_o,_al_u865_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(0*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)))"),
    //.LUTF1("(~(A)*~(C)*~(B)*D*~(0)+A*~(C)*~(B)*D*~(0)+~(A)*C*~(B)*D*~(0)+~(A)*~(C)*B*D*~(0)+A*~(C)*B*D*~(0)+~(A)*C*B*D*~(0)+~(A)*~(C)*~(B)*~(D)*0+A*~(C)*~(B)*~(D)*0+~(A)*C*~(B)*~(D)*0+~(A)*~(C)*B*~(D)*0+A*~(C)*B*~(D)*0+~(A)*C*B*~(D)*0+~(A)*~(C)*~(B)*D*0+A*~(C)*~(B)*D*0+~(A)*C*~(B)*D*0+A*C*~(B)*D*0+~(A)*~(C)*B*D*0+A*~(C)*B*D*0)"),
    //.LUTG0("~(~A*~(1*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)))"),
    //.LUTG1("(~(A)*~(C)*~(B)*D*~(1)+A*~(C)*~(B)*D*~(1)+~(A)*C*~(B)*D*~(1)+~(A)*~(C)*B*D*~(1)+A*~(C)*B*D*~(1)+~(A)*C*B*D*~(1)+~(A)*~(C)*~(B)*~(D)*1+A*~(C)*~(B)*~(D)*1+~(A)*C*~(B)*~(D)*1+~(A)*~(C)*B*~(D)*1+A*~(C)*B*~(D)*1+~(A)*C*B*~(D)*1+~(A)*~(C)*~(B)*D*1+A*~(C)*~(B)*D*1+~(A)*C*~(B)*D*1+A*C*~(B)*D*1+~(A)*~(C)*B*D*1+A*~(C)*B*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b0101111100000000),
    .INIT_LUTG0(16'b1110111011111010),
    .INIT_LUTG1(16'b0011111101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u853|picorv32_core/reg14_b20  (
    .a({_al_u826_o,_al_u853_o}),
    .b({_al_u828_o,\picorv32_core/n433 [20]}),
    .c({_al_u827_o,\picorv32_core/n434 [20]}),
    .clk(clk_pad),
    .d({\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/instr_sub }),
    .e({\picorv32_core/pcpi_rs2$20$ ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u853_o,open_n19211}),
    .q({open_n19215,\picorv32_core/alu_out_q [20]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .INIT_LUT0(16'b0111011100000000),
    .INIT_LUT1(16'b0011111101110111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u857 (
    .a({_al_u826_o,_al_u826_o}),
    .b({_al_u827_o,_al_u827_o}),
    .c({_al_u828_o,_al_u828_o}),
    .d({\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs1$22$ }),
    .mi({open_n19228,\picorv32_core/pcpi_rs2$22$ }),
    .fx({open_n19233,_al_u857_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(0*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)))"),
    //.LUTF1("~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+~D*~B*C*A+D*~B*C*A+~D*B*C*A"),
    //.LUTG0("~(~D*~(1*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)))"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+~D*~B*C*A+D*~B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b1111111111001010),
    .INIT_LUTG1(16'b0111001101111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u859|picorv32_core/reg14_b23  (
    .a({_al_u828_o,\picorv32_core/n434 [23]}),
    .b({_al_u827_o,\picorv32_core/n433 [23]}),
    .c({\picorv32_core/pcpi_rs2$23$ ,\picorv32_core/instr_sub }),
    .clk(clk_pad),
    .d({_al_u826_o,_al_u859_o}),
    .e({\picorv32_core/pcpi_rs1$23$ ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u859_o,open_n19252}),
    .q({open_n19256,\picorv32_core/alu_out_q [23]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(0*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)))"),
    //.LUTF1("~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D"),
    //.LUTG0("~(~A*~(1*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)))"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b0101111100000000),
    .INIT_LUTG0(16'b1110111011111010),
    .INIT_LUTG1(16'b0011111101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u861|picorv32_core/reg14_b24  (
    .a({_al_u826_o,_al_u861_o}),
    .b({_al_u828_o,\picorv32_core/n433 [24]}),
    .c({_al_u827_o,\picorv32_core/n434 [24]}),
    .clk(clk_pad),
    .d({\picorv32_core/pcpi_rs2$24$ ,\picorv32_core/instr_sub }),
    .e({\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u861_o,open_n19273}),
    .q({open_n19277,\picorv32_core/alu_out_q [24]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .INIT_LUT0(16'b0111011100000000),
    .INIT_LUT1(16'b0011111101110111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u863 (
    .a({_al_u826_o,_al_u826_o}),
    .b({_al_u827_o,_al_u827_o}),
    .c({_al_u828_o,_al_u828_o}),
    .d({\picorv32_core/pcpi_rs1$25$ ,\picorv32_core/pcpi_rs1$25$ }),
    .mi({open_n19290,\picorv32_core/pcpi_rs2$25$ }),
    .fx({open_n19295,_al_u863_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(0*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)))"),
    //.LUTF1("~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D"),
    //.LUTG0("~(~A*~(1*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)))"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b0101111100000000),
    .INIT_LUTG0(16'b1110111011111010),
    .INIT_LUTG1(16'b0011111101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u867|picorv32_core/reg14_b27  (
    .a({_al_u826_o,_al_u867_o}),
    .b({_al_u828_o,\picorv32_core/n433 [27]}),
    .c({_al_u827_o,\picorv32_core/n434 [27]}),
    .clk(clk_pad),
    .d({\picorv32_core/pcpi_rs2$27$ ,\picorv32_core/instr_sub }),
    .e({\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u867_o,open_n19314}),
    .q({open_n19318,\picorv32_core/alu_out_q [27]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(0*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)))"),
    //.LUTF1("~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+~D*~B*C*A+D*~B*C*A+~D*B*C*A"),
    //.LUTG0("~(~D*~(1*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)))"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+~D*~B*C*A+D*~B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b1111111111001010),
    .INIT_LUTG1(16'b0111001101111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u869|picorv32_core/reg14_b28  (
    .a({_al_u828_o,\picorv32_core/n434 [28]}),
    .b({_al_u827_o,\picorv32_core/n433 [28]}),
    .c({\picorv32_core/pcpi_rs2$28$ ,\picorv32_core/instr_sub }),
    .clk(clk_pad),
    .d({_al_u826_o,_al_u869_o}),
    .e({\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u869_o,open_n19335}),
    .q({open_n19339,\picorv32_core/alu_out_q [28]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .INIT_LUT0(16'b0111011100000000),
    .INIT_LUT1(16'b0011111101110111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u871 (
    .a({_al_u826_o,_al_u826_o}),
    .b({_al_u827_o,_al_u827_o}),
    .c({_al_u828_o,_al_u828_o}),
    .d({\picorv32_core/pcpi_rs1$29$ ,\picorv32_core/pcpi_rs1$29$ }),
    .mi({open_n19352,\picorv32_core/pcpi_rs2$29$ }),
    .fx({open_n19357,_al_u871_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(0*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)))"),
    //.LUTF1("(~(A)*~(C)*~(B)*D*~(0)+A*~(C)*~(B)*D*~(0)+~(A)*C*~(B)*D*~(0)+~(A)*~(C)*B*D*~(0)+A*~(C)*B*D*~(0)+~(A)*C*B*D*~(0)+~(A)*~(C)*~(B)*~(D)*0+A*~(C)*~(B)*~(D)*0+~(A)*C*~(B)*~(D)*0+~(A)*~(C)*B*~(D)*0+A*~(C)*B*~(D)*0+~(A)*C*B*~(D)*0+~(A)*~(C)*~(B)*D*0+A*~(C)*~(B)*D*0+~(A)*C*~(B)*D*0+A*C*~(B)*D*0+~(A)*~(C)*B*D*0+A*~(C)*B*D*0)"),
    //.LUTG0("~(~A*~(1*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)))"),
    //.LUTG1("(~(A)*~(C)*~(B)*D*~(1)+A*~(C)*~(B)*D*~(1)+~(A)*C*~(B)*D*~(1)+~(A)*~(C)*B*D*~(1)+A*~(C)*B*D*~(1)+~(A)*C*B*D*~(1)+~(A)*~(C)*~(B)*~(D)*1+A*~(C)*~(B)*~(D)*1+~(A)*C*~(B)*~(D)*1+~(A)*~(C)*B*~(D)*1+A*~(C)*B*~(D)*1+~(A)*C*B*~(D)*1+~(A)*~(C)*~(B)*D*1+A*~(C)*~(B)*D*1+~(A)*C*~(B)*D*1+A*C*~(B)*D*1+~(A)*~(C)*B*D*1+A*~(C)*B*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b0101111100000000),
    .INIT_LUTG0(16'b1110111011111010),
    .INIT_LUTG1(16'b0011111101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u875|picorv32_core/reg14_b30  (
    .a({_al_u826_o,_al_u875_o}),
    .b({_al_u828_o,\picorv32_core/n433 [30]}),
    .c({_al_u827_o,\picorv32_core/n434 [30]}),
    .clk(clk_pad),
    .d({\picorv32_core/pcpi_rs1$30$ ,\picorv32_core/instr_sub }),
    .e({\picorv32_core/pcpi_rs2$30$ ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u875_o,open_n19376}),
    .q({open_n19380,\picorv32_core/alu_out_q [30]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(0*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)))"),
    //.LUTF1("~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+~D*~B*C*A+D*~B*C*A+~D*B*C*A"),
    //.LUTG0("~(~D*~(1*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)))"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+~D*~B*C*A+D*~B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b1111111111001010),
    .INIT_LUTG1(16'b0111001101111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u877|picorv32_core/reg14_b31  (
    .a({_al_u828_o,\picorv32_core/n434 [31]}),
    .b({_al_u827_o,\picorv32_core/n433 [31]}),
    .c({\picorv32_core/pcpi_rs2$31$ ,\picorv32_core/instr_sub }),
    .clk(clk_pad),
    .d({_al_u826_o,_al_u877_o}),
    .e({\picorv32_core/pcpi_rs1$31$ ,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .f({_al_u877_o,open_n19397}),
    .q({open_n19401,\picorv32_core/alu_out_q [31]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(C)*~(B)*~(D)*A*~(1)+C*~(B)*~(D)*A*~(1)+~(C)*B*~(D)*A*~(1)+~(C)*~(B)*D*A*~(1)+C*~(B)*D*A*~(1)+~(C)*B*D*A*~(1)+~(C)*~(B)*~(D)*~(A)*1+C*~(B)*~(D)*~(A)*1+~(C)*B*~(D)*~(A)*1+~(C)*~(B)*D*~(A)*1+C*~(B)*D*~(A)*1+~(C)*B*D*~(A)*1+~(C)*~(B)*~(D)*A*1+C*~(B)*~(D)*A*1+~(C)*B*~(D)*A*1+C*B*~(D)*A*1+~(C)*~(B)*D*A*1+C*~(B)*D*A*1)"),
    .INIT_LUT0(16'b0111011100000000),
    .INIT_LUT1(16'b0011011110111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u887 (
    .a({\picorv32_core/pcpi_rs1$8$ ,_al_u826_o}),
    .b({_al_u827_o,_al_u827_o}),
    .c({_al_u826_o,_al_u828_o}),
    .d({_al_u828_o,\picorv32_core/pcpi_rs1$8$ }),
    .mi({open_n19414,\picorv32_core/pcpi_rs2$8$ }),
    .fx({open_n19419,_al_u887_o}));
  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~A)"),
    //.LUT1("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111101011111010),
    .INIT_LUT1(16'b0100010101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u894|uart/reg6_b0  (
    .a({\uart/uart_idr [0],\uart/mux51_b0_sel_is_3_o }),
    .b({\picorv32_core/pcpi_rs1$2$ ,open_n19422}),
    .c({_al_u700_o_placeOpt_1,\uart/uart_status_rx_clr }),
    .ce(\uart/mux51_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\picorv32_core/n30 [0],open_n19423}),
    .mi({open_n19434,\uart/uart_idr_t [0]}),
    .sr(resetn_placeOpt_8),
    .f({_al_u894_o,\picorv32_core/n524$4$_en }),
    .q({open_n19438,\uart/uart_idr [0]}));  // ../src/uart.v(263)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D"),
    //.LUTG1("~B*~C*~A*~D+B*~C*~A*~D+~B*~C*~A*D+B*~C*~A*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010101010101),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0111011101110111),
    .INIT_LUTG1(16'b0000010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u896|picorv32_core/reg11_b2  (
    .a({\picorv32_core/is_sb_sh_sw ,_al_u906_o}),
    .b({open_n19439,_al_u803_o}),
    .c({\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ,open_n19440}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .e({_al_u803_o,\picorv32_core/mem_rdata_q [22]}),
    .f({_al_u896_o,open_n19458}),
    .q({open_n19462,\picorv32_core/decoded_imm [2]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~(~C*~B))*~(0*A))"),
    //.LUT1("(~(B*~(~C*~D))*~(1*A))"),
    .INIT_LUT0(16'b0000001111111111),
    .INIT_LUT1(16'b0001000100010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u904 (
    .a({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .b({\picorv32_core/mem_rdata_q [10],\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .c({\picorv32_core/is_sb_sh_sw ,\picorv32_core/is_sb_sh_sw }),
    .d({\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ,\picorv32_core/mem_rdata_q [10]}),
    .mi({open_n19475,\picorv32_core/decoded_imm_uj [3]}),
    .fx({open_n19480,_al_u904_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~(~C*~B))*~(0*A))"),
    //.LUT1("(~(B*~(~C*~D))*~(1*A))"),
    .INIT_LUT0(16'b0000001111111111),
    .INIT_LUT1(16'b0001000100010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u906 (
    .a({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .b({\picorv32_core/mem_rdata_q [9],\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .c({\picorv32_core/is_sb_sh_sw ,\picorv32_core/is_sb_sh_sw }),
    .d({\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ,\picorv32_core/mem_rdata_q [9]}),
    .mi({open_n19495,\picorv32_core/decoded_imm_uj [2]}),
    .fx({open_n19500,_al_u906_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~A*~(C*B))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0001010100010101),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0001010100010101),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u908|_al_u909  (
    .a({open_n19503,_al_u908_o}),
    .b({open_n19504,\picorv32_core/instr_jal }),
    .c({\picorv32_core/mem_rdata_q [31],\picorv32_core/decoded_imm_uj [20]}),
    .d({_al_u896_o,open_n19507}),
    .f({_al_u908_o,_al_u909_o}));
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(A*~(~C*B)))"),
    //.LUT1("(~(A*D)*~(B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010001011111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u930|picorv32_core/reg11_b11  (
    .a({\picorv32_core/mem_rdata_q [7],\picorv32_core/mem_rdata_q [31]}),
    .b({\picorv32_core/decoded_imm_uj [11],_al_u803_o}),
    .c({\picorv32_core/instr_jal ,\picorv32_core/is_sb_sh_sw }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ,_al_u930_o}),
    .f({_al_u930_o,open_n19543}),
    .q({open_n19547,\picorv32_core/decoded_imm [11]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(B*D)"),
    //.LUT1("(~A*C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110000000000),
    .INIT_LUT1(16'b0000000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u960|picorv32_core/instr_sw_reg  (
    .a({\picorv32_core/mem_rdata_q [14],open_n19548}),
    .b({open_n19549,\picorv32_core/is_sb_sh_sw }),
    .c({\picorv32_core/mem_rdata_q [13],open_n19550}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [12],\picorv32_core/n289_lutinv }),
    .f({\picorv32_core/n289_lutinv ,open_n19564}),
    .q({open_n19568,\picorv32_core/instr_sw }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)"),
    //.LUT1("(D*B)"),
    .INIT_LUT0(16'b1100110010101010),
    .INIT_LUT1(16'b1100110000000000),
    .MODE("LOGIC"))
    \_al_u976|_al_u1226  (
    .a({open_n19569,\uart/n49 [1]}),
    .b({\picorv32_core/n304_lutinv ,\uart/uart_smp_rx [1]}),
    .d({\picorv32_core/is_alu_reg_reg ,rxd_pad}),
    .f({_al_u976_o,\uart/n50 [1]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~C*D))"),
    //.LUT1("(~D*~B*~C)"),
    .INIT_LUT0(16'b1010000010101010),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"))
    \_al_u979|_al_u1555  (
    .a({open_n19592,_al_u1554_o}),
    .b({\picorv32_core/cpu_state [1],open_n19593}),
    .c({\picorv32_core/cpu_state [0],_al_u1551_o}),
    .d({\picorv32_core/cpu_state [2],\picorv32_core/n523_lutinv }),
    .f({_al_u979_o,_al_u1555_o}));
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    //.LUTF1("(~D*~C)"),
    //.LUTG0("0"),
    //.LUTG1("(~D*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u980|picorv32_core/reg22_b5  (
    .b({open_n19616,\picorv32_core/sel39_b0_sel_is_3_o }),
    .c({1'b0,resetn_placeOpt_8}),
    .clk(clk_pad),
    .d({\picorv32_core/cpu_state [5],open_n19618}),
    .e({open_n19619,\picorv32_core/instr_jal }),
    .sr(\picorv32_core/mux164_b0_sel_is_0_o ),
    .f({_al_u980_o,open_n19634}),
    .q({open_n19638,\picorv32_core/cpu_state [5]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~0*A*~C*B*D)"),
    //.LUT1("(~1*A*~C*B*D)"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u981 (
    .a({\picorv32_core/cpu_state [6],\picorv32_core/cpu_state [6]}),
    .b({_al_u980_o,_al_u980_o}),
    .c({\picorv32_core/cpu_state [3],\picorv32_core/cpu_state [3]}),
    .d({_al_u979_o,_al_u979_o}),
    .mi({open_n19651,\picorv32_core/cpu_state [7]}),
    .fx({open_n19656,\picorv32_core/n663 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u982|_al_u1152  (
    .b({open_n19661,_al_u979_o}),
    .c({\picorv32_core/cpu_state [3],\picorv32_core/cpu_state [3]}),
    .d({_al_u979_o,_al_u1147_o}),
    .f({_al_u982_o,\picorv32_core/n666_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~0*B*~C*~D*A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~1*B*~C*~D*A)"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u992|_al_u974  (
    .a({_al_u973_o,_al_u973_o}),
    .b({\picorv32_core/mem_rdata_q [30],\picorv32_core/mem_rdata_q [28]}),
    .c({\picorv32_core/mem_rdata_q [29],\picorv32_core/mem_rdata_q [29]}),
    .d({\picorv32_core/mem_rdata_q [28],\picorv32_core/mem_rdata_q [30]}),
    .e({\picorv32_core/mem_rdata_q [31],\picorv32_core/mem_rdata_q [31]}),
    .f({\picorv32_core/n308_lutinv ,\picorv32_core/n304_lutinv }));
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*B*A)"),
    //.LUTF1("0"),
    //.LUTG0("(~1*~D*~C*B*A)"),
    //.LUTG1("~C*B*~D*A+C*B*~D*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u993|picorv32_core/instr_sub_reg  (
    .a({\picorv32_core/mem_rdata_q [14],\picorv32_core/n308_lutinv }),
    .b({\picorv32_core/mem_rdata_q [12],\picorv32_core/is_alu_reg_reg }),
    .c({open_n19704,\picorv32_core/mem_rdata_q [12]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [13],\picorv32_core/mem_rdata_q [13]}),
    .e({\picorv32_core/n308_lutinv ,\picorv32_core/mem_rdata_q [14]}),
    .sr(resetn_placeOpt_16),
    .f({\picorv32_core/n345 ,open_n19719}),
    .q({open_n19723,\picorv32_core/instr_sub }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*~(A)*~(B)+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*~(B)+~((D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C))*A*B+(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)*A*B)"),
    //.LUT1("~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*~(A)*~(B)+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*~(B)+~((D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C))*A*B+(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)*A*B)"),
    .INIT_LUT0(16'b0111010001110111),
    .INIT_LUT1(16'b0100010001000111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u999 (
    .a({\picorv32_core/n450 [9],\picorv32_core/n450 [9]}),
    .b({\picorv32_core/latched_branch ,\picorv32_core/latched_branch }),
    .c({\picorv32_core/latched_stalu ,\picorv32_core/latched_stalu }),
    .d({\picorv32_core/reg_out [9],\picorv32_core/reg_out [9]}),
    .mi({open_n19736,\picorv32_core/alu_out_q [9]}),
    .fx({open_n19741,_al_u999_o}));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0004"),
    //.WID("0x0004"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0185F7C7100007078BF7C71000C68044FB0F00070700FE070707101131800000),
    .INIT_01(256'h44FEFB278047FEFE97272722FEA0222426CE80540000FD3F00FC00FDA82ED471),
    .INIT_02(256'h44003C3F053708C680544745272726FEA80000972627C7FDFEA8262A2C2ED680),
    .INIT_03(256'hC680540085C7FF8B4785C7FF0F8347062487472287472087372E87370700DE80),
    .INIT_04(256'h2785F7FD3D0585F72785F7FE3F0F872785F7FE3D0524272C2ED4710140353508),
    .INIT_05(256'h2702350097272702350FFE3D0F872785F7FE350F8727FE9727278B27FE3F85F7),
    .INIT_06(256'h566900FE69672724FCA02407FE00FE1035060407070724DC716150F8FDFEFE07),
    .INIT_07(256'h307A006D206D70000A7461632E00742072392E00383047617220676E29203228),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000031292843),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \mem_hi/inst_1024x8_sub_000000_000  (
    .addra({mem_la_addr[11:2],3'b111}),
    .clka(clk_pad),
    .dia({open_n19813,mem_la_wdata[31:24]}),
    .rsta(resetn_placeOpt_15),
    .wea(n13),
    .doa({open_n19827,memory_out[31:24]}));
  // address_offset=0;data_offset=0;depth=1024;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0005"),
    //.WID("0x0005"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h32F707D1B72300E5F707F1B7004105018593830001230300F4AA2202EF133700),
    .INIT_01(256'h3E8344E707368303C444F4FD83C4B4A4000145B2F583833E83231383A4000682),
    .INIT_02(256'hB229134019132241453EF744C4F4858381638384C407BA038304C4B4A4007905),
    .INIT_03(256'h4121F20DC7BA13F41DC7BA1393F404F43745F48741F44736F40732F4AA223941),
    .INIT_04(256'h21F7A1838031F74425F7A1833E934491F7E18340F4C4B4A40006822201293522),
    .INIT_05(256'h19133E8384C43D133E93833E9344C1F7C1833E93449123C4C4B9C4A523F5F784),
    .INIT_06(256'h630DF1E39384F4858304F485832303B70498130004048006822201E3830323C4),
    .INIT_07(256'h652020666F2044000D2E6873770D7069203241294E34646B53206E2049495233),
    .INIT_08(256'h00000000000000000000000000000000000000000000000000002E2E20474378),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \mem_lo/inst_1024x8_sub_000000_000  (
    .addra({mem_la_addr[11:2],3'b111}),
    .clka(clk_pad),
    .dia({open_n19859,mem_la_wdata[7:0]}),
    .rsta(resetn_placeOpt_15),
    .wea(n7),
    .doa({open_n19873,memory_out[7:0]}));
  // address_offset=0;data_offset=0;depth=1024;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0006"),
    //.WID("0x0006"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h413E93830007F1B78993830001228272E5F707F1B7E7F4C1B7A3000120010000),
    .INIT_01(256'h72C4F98323038444BA03832344252323232282220107C48507E417C419232279),
    .INIT_02(256'h2201C00113800006823285E3830323C429F707B6838303C4C405232323232282),
    .INIT_03(256'h068262013E8304BD833E8304F79183232393B72393B72393B72393B7A3800682),
    .INIT_04(256'h833E938411133E93833E93441DF7C1833E9344811323832323227941B2213100),
    .INIT_05(256'h83007907BA0383005DF7444DF7A1833E9344F9F7E183F4BA8303BD83048D3E93),
    .INIT_06(256'h525000E7F7E10323843123A3F4E7F4000D2350E1B7A323223945B2F784C4F485),
    .INIT_07(256'h2069786F79656D000D656E637700726C6531720A3832456F616E6E7541433320),
    .INIT_08(256'h000000000000000000000000000000000000000000000000000000002E552047),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \mem_mh/inst_1024x8_sub_000000_000  (
    .addra({mem_la_addr[11:2],3'b111}),
    .clka(clk_pad),
    .dia({open_n19905,mem_la_wdata[23:16]}),
    .rsta(resetn_placeOpt_15),
    .wea(n11),
    .doa({open_n19919,memory_out[23:16]}));
  // address_offset=0;data_offset=0;depth=1024;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0007"),
    //.WID("0x0007"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h440F0007078010DB0F000707081161008BF7C71000804710FE87CE9000011100),
    .INIT_01(256'h8527FE0000972627FEFEFE1727FEFEFE10116150F3C72785C72E8727FC18D680),
    .INIT_02(256'h4037053B3F05C4116185FCFDFEFE07274704C7FDFE00972727FEFCFCFC187161),
    .INIT_03(256'h11615035FE9707FC3DFE9707F7FCFEFE4446FE9342FE5337FC1333FC87DC7101),
    .INIT_04(256'h370F87273F3F0FFE370F872785F7FE370F87273EFEFDFCFC18D68044004545C4),
    .INIT_05(256'h3B0585C7FEFE330585F72785F7FE350F872785F7FE3F22FEFDE7FEA8263D0FFD),
    .INIT_06(256'h6F0AB7D687FCFC0727FCFE0747804707FCC30710FEFC00DE80540041272726FE),
    .INIT_07(256'h3A733072726D75000A6E696F770A6F615330700D47532852706F6972534D5632),
    .INIT_08(256'h00000000000000000000000000000000000000000000000000003030364E3A00),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("INV"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \mem_ml/inst_1024x8_sub_000000_000  (
    .addra({mem_la_addr[11:2],3'b111}),
    .clka(clk_pad),
    .dia({open_n19951,mem_la_wdata[15:8]}),
    .rsta(resetn_placeOpt_2),
    .wea(n9),
    .doa({open_n19965,memory_out[15:8]}));
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P11"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("RESET"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("1"),
    .OUTRSTMUX("INV"),
    .OUTSCLKMUX("CLK"),
    .SRMODE("ASYNC"),
    .TSMUX("0"))
    out_byte_en_reg_DO (
    .ce(1'b1),
    .do({open_n19975,open_n19976,open_n19977,n16}),
    .osclk(clk_pad),
    .rst(resetn_placeOpt_4),
    .opad(out_byte_en));  // ../src/top.v(128)
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u0|picorv32_core/add0/ucin  (
    .a({\picorv32_core/next_pc [2],1'b0}),
    .b({\picorv32_core/mem_la_firstword_xfer ,open_n19989}),
    .f({\picorv32_core/n30 [0],open_n20009}),
    .fco(\picorv32_core/add0/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u10|picorv32_core/add0/u9  (
    .a({\picorv32_core/next_pc [12],1'b0}),
    .b({1'b0,\picorv32_core/next_pc [11]}),
    .fci(\picorv32_core/add0/c9 ),
    .f(\picorv32_core/n30 [10:9]),
    .fco(\picorv32_core/add0/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u12|picorv32_core/add0/u11  (
    .a({1'b0,\picorv32_core/next_pc [13]}),
    .b({\picorv32_core/next_pc [14],1'b0}),
    .fci(\picorv32_core/add0/c11 ),
    .f(\picorv32_core/n30 [12:11]),
    .fco(\picorv32_core/add0/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u14|picorv32_core/add0/u13  (
    .a(2'b00),
    .b(\picorv32_core/next_pc [16:15]),
    .fci(\picorv32_core/add0/c13 ),
    .f(\picorv32_core/n30 [14:13]),
    .fco(\picorv32_core/add0/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u16|picorv32_core/add0/u15  (
    .a({\picorv32_core/next_pc [18],1'b0}),
    .b({1'b0,\picorv32_core/next_pc [17]}),
    .fci(\picorv32_core/add0/c15 ),
    .f(\picorv32_core/n30 [16:15]),
    .fco(\picorv32_core/add0/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u18|picorv32_core/add0/u17  (
    .a(\picorv32_core/next_pc [20:19]),
    .b(2'b00),
    .fci(\picorv32_core/add0/c17 ),
    .f(\picorv32_core/n30 [18:17]),
    .fco(\picorv32_core/add0/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u20|picorv32_core/add0/u19  (
    .a({\picorv32_core/next_pc [22],1'b0}),
    .b({1'b0,\picorv32_core/next_pc [21]}),
    .fci(\picorv32_core/add0/c19 ),
    .f(\picorv32_core/n30 [20:19]),
    .fco(\picorv32_core/add0/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u22|picorv32_core/add0/u21  (
    .a(2'b00),
    .b(\picorv32_core/next_pc [24:23]),
    .fci(\picorv32_core/add0/c21 ),
    .f(\picorv32_core/n30 [22:21]),
    .fco(\picorv32_core/add0/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u24|picorv32_core/add0/u23  (
    .a(\picorv32_core/next_pc [26:25]),
    .b(2'b00),
    .fci(\picorv32_core/add0/c23 ),
    .f(\picorv32_core/n30 [24:23]),
    .fco(\picorv32_core/add0/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u26|picorv32_core/add0/u25  (
    .a({\picorv32_core/next_pc [28],1'b0}),
    .b({1'b0,\picorv32_core/next_pc [27]}),
    .fci(\picorv32_core/add0/c25 ),
    .f(\picorv32_core/n30 [26:25]),
    .fco(\picorv32_core/add0/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u28|picorv32_core/add0/u27  (
    .a(\picorv32_core/next_pc [30:29]),
    .b(2'b00),
    .fci(\picorv32_core/add0/c27 ),
    .f(\picorv32_core/n30 [28:27]),
    .fco(\picorv32_core/add0/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u29_al_u2574  (
    .a({open_n20234,\picorv32_core/next_pc [31]}),
    .b({open_n20235,1'b0}),
    .fci(\picorv32_core/add0/c29 ),
    .f({open_n20254,\picorv32_core/n30 [29]}));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u2|picorv32_core/add0/u1  (
    .a({1'b0,\picorv32_core/next_pc [3]}),
    .b({\picorv32_core/next_pc [4],1'b0}),
    .fci(\picorv32_core/add0/c1 ),
    .f(\picorv32_core/n30 [2:1]),
    .fco(\picorv32_core/add0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u4|picorv32_core/add0/u3  (
    .a({1'b0,\picorv32_core/next_pc [5]}),
    .b({\picorv32_core/next_pc [6],1'b0}),
    .fci(\picorv32_core/add0/c3 ),
    .f(\picorv32_core/n30 [4:3]),
    .fco(\picorv32_core/add0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u6|picorv32_core/add0/u5  (
    .a(2'b00),
    .b(\picorv32_core/next_pc [8:7]),
    .fci(\picorv32_core/add0/c5 ),
    .f(\picorv32_core/n30 [6:5]),
    .fco(\picorv32_core/add0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add0/u0|picorv32_core/add0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add0/u8|picorv32_core/add0/u7  (
    .a(2'b00),
    .b(\picorv32_core/next_pc [10:9]),
    .fci(\picorv32_core/add0/c7 ),
    .f(\picorv32_core/n30 [8:7]),
    .fco(\picorv32_core/add0/c9 ));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add1/ucin_al_u2529"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add1/u11_al_u2532  (
    .a({\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/pcpi_rs1$11$ }),
    .b({\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$12$ }),
    .c(2'b00),
    .d({\picorv32_core/pcpi_rs2$13$ ,\picorv32_core/pcpi_rs2$11$ }),
    .e({\picorv32_core/pcpi_rs2$14$ ,\picorv32_core/pcpi_rs2$12$ }),
    .fci(\picorv32_core/add1/c11 ),
    .f({\picorv32_core/n434 [13],\picorv32_core/n434 [11]}),
    .fco(\picorv32_core/add1/c15 ),
    .fx({\picorv32_core/n434 [14],\picorv32_core/n434 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add1/ucin_al_u2529"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add1/u15_al_u2533  (
    .a({\picorv32_core/pcpi_rs1$17$ ,\picorv32_core/pcpi_rs1$15$ }),
    .b({\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$16$ }),
    .c(2'b00),
    .d({\picorv32_core/pcpi_rs2$17$ ,\picorv32_core/pcpi_rs2$15$ }),
    .e({\picorv32_core/pcpi_rs2$18$ ,\picorv32_core/pcpi_rs2$16$ }),
    .fci(\picorv32_core/add1/c15 ),
    .f({\picorv32_core/n434 [17],\picorv32_core/n434 [15]}),
    .fco(\picorv32_core/add1/c19 ),
    .fx({\picorv32_core/n434 [18],\picorv32_core/n434 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add1/ucin_al_u2529"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add1/u19_al_u2534  (
    .a({\picorv32_core/pcpi_rs1$21$ ,\picorv32_core/pcpi_rs1$19$ }),
    .b({\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs1$20$ }),
    .c(2'b00),
    .d({\picorv32_core/pcpi_rs2$21$ ,\picorv32_core/pcpi_rs2$19$ }),
    .e({\picorv32_core/pcpi_rs2$22$ ,\picorv32_core/pcpi_rs2$20$ }),
    .fci(\picorv32_core/add1/c19 ),
    .f({\picorv32_core/n434 [21],\picorv32_core/n434 [19]}),
    .fco(\picorv32_core/add1/c23 ),
    .fx({\picorv32_core/n434 [22],\picorv32_core/n434 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add1/ucin_al_u2529"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add1/u23_al_u2535  (
    .a({\picorv32_core/pcpi_rs1$25$ ,\picorv32_core/pcpi_rs1$23$ }),
    .b({\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$24$ }),
    .c(2'b00),
    .d({\picorv32_core/pcpi_rs2$25$ ,\picorv32_core/pcpi_rs2$23$ }),
    .e({\picorv32_core/pcpi_rs2$26$ ,\picorv32_core/pcpi_rs2$24$ }),
    .fci(\picorv32_core/add1/c23 ),
    .f({\picorv32_core/n434 [25],\picorv32_core/n434 [23]}),
    .fco(\picorv32_core/add1/c27 ),
    .fx({\picorv32_core/n434 [26],\picorv32_core/n434 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add1/ucin_al_u2529"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add1/u27_al_u2536  (
    .a({\picorv32_core/pcpi_rs1$29$ ,\picorv32_core/pcpi_rs1$27$ }),
    .b({\picorv32_core/pcpi_rs1$30$ ,\picorv32_core/pcpi_rs1$28$ }),
    .c(2'b00),
    .d({\picorv32_core/pcpi_rs2$29$ ,\picorv32_core/pcpi_rs2$27$ }),
    .e({\picorv32_core/pcpi_rs2$30$ ,\picorv32_core/pcpi_rs2$28$ }),
    .fci(\picorv32_core/add1/c27 ),
    .f({\picorv32_core/n434 [29],\picorv32_core/n434 [27]}),
    .fco(\picorv32_core/add1/c31 ),
    .fx({\picorv32_core/n434 [30],\picorv32_core/n434 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add1/ucin_al_u2529"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add1/u31_al_u2537  (
    .a({open_n20438,\picorv32_core/pcpi_rs1$31$ }),
    .c(2'b00),
    .d({open_n20443,\picorv32_core/pcpi_rs2$31$ }),
    .fci(\picorv32_core/add1/c31 ),
    .f({open_n20460,\picorv32_core/n434 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add1/ucin_al_u2529"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add1/u3_al_u2530  (
    .a({\picorv32_core/pcpi_rs1$5$ ,\picorv32_core/pcpi_rs1$3$ }),
    .b({\picorv32_core/pcpi_rs1$6$ ,\picorv32_core/pcpi_rs1$4$ }),
    .c(2'b00),
    .d({mem_la_wdata[5],mem_la_wdata[3]}),
    .e({mem_la_wdata[6],mem_la_wdata[4]}),
    .fci(\picorv32_core/add1/c3 ),
    .f({\picorv32_core/n434 [5],\picorv32_core/n434 [3]}),
    .fco(\picorv32_core/add1/c7 ),
    .fx({\picorv32_core/n434 [6],\picorv32_core/n434 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add1/ucin_al_u2529"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add1/u7_al_u2531  (
    .a({\picorv32_core/pcpi_rs1$9$ ,\picorv32_core/pcpi_rs1$7$ }),
    .b({\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$8$ }),
    .c(2'b00),
    .d({\picorv32_core/pcpi_rs2$9$ ,mem_la_wdata[7]}),
    .e({\picorv32_core/pcpi_rs2$10$ ,\picorv32_core/pcpi_rs2$8$ }),
    .fci(\picorv32_core/add1/c7 ),
    .f({\picorv32_core/n434 [9],\picorv32_core/n434 [7]}),
    .fco(\picorv32_core/add1/c11 ),
    .fx({\picorv32_core/n434 [10],\picorv32_core/n434 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add1/ucin_al_u2529"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \picorv32_core/add1/ucin_al_u2529  (
    .a({\picorv32_core/pcpi_rs1$1$ ,1'b0}),
    .b({\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$0$ }),
    .c(2'b00),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({mem_la_wdata[1],1'b1}),
    .e({mem_la_wdata[2],mem_la_wdata[0]}),
    .mi(mem_la_wdata[2:1]),
    .sr(resetn),
    .f({\picorv32_core/n434 [1],open_n20514}),
    .fco(\picorv32_core/add1/c3 ),
    .fx({\picorv32_core/n434 [2],\picorv32_core/n434 [0]}),
    .q(\uart/uart_bsrr [2:1]));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add2/ucin_al_u2538"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add2/u11_al_u2541  (
    .a({\picorv32_core/reg_pc [13],\picorv32_core/reg_pc [11]}),
    .b({\picorv32_core/reg_pc [14],\picorv32_core/reg_pc [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add2/c11 ),
    .f({\picorv32_core/n450 [13],\picorv32_core/n450 [11]}),
    .fco(\picorv32_core/add2/c15 ),
    .fx({\picorv32_core/n450 [14],\picorv32_core/n450 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add2/ucin_al_u2538"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add2/u15_al_u2542  (
    .a({\picorv32_core/reg_pc [17],\picorv32_core/reg_pc [15]}),
    .b({\picorv32_core/reg_pc [18],\picorv32_core/reg_pc [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add2/c15 ),
    .f({\picorv32_core/n450 [17],\picorv32_core/n450 [15]}),
    .fco(\picorv32_core/add2/c19 ),
    .fx({\picorv32_core/n450 [18],\picorv32_core/n450 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add2/ucin_al_u2538"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add2/u19_al_u2543  (
    .a({\picorv32_core/reg_pc [21],\picorv32_core/reg_pc [19]}),
    .b({\picorv32_core/reg_pc [22],\picorv32_core/reg_pc [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add2/c19 ),
    .f({\picorv32_core/n450 [21],\picorv32_core/n450 [19]}),
    .fco(\picorv32_core/add2/c23 ),
    .fx({\picorv32_core/n450 [22],\picorv32_core/n450 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add2/ucin_al_u2538"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add2/u23_al_u2544  (
    .a({\picorv32_core/reg_pc [25],\picorv32_core/reg_pc [23]}),
    .b({\picorv32_core/reg_pc [26],\picorv32_core/reg_pc [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add2/c23 ),
    .f({\picorv32_core/n450 [25],\picorv32_core/n450 [23]}),
    .fco(\picorv32_core/add2/c27 ),
    .fx({\picorv32_core/n450 [26],\picorv32_core/n450 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add2/ucin_al_u2538"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add2/u27_al_u2545  (
    .a({\picorv32_core/reg_pc [29],\picorv32_core/reg_pc [27]}),
    .b({\picorv32_core/reg_pc [30],\picorv32_core/reg_pc [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add2/c27 ),
    .f({\picorv32_core/n450 [29],\picorv32_core/n450 [27]}),
    .fco(\picorv32_core/add2/c31 ),
    .fx({\picorv32_core/n450 [30],\picorv32_core/n450 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add2/ucin_al_u2538"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add2/u31_al_u2546  (
    .a({open_n20605,\picorv32_core/reg_pc [31]}),
    .c(2'b00),
    .d({open_n20610,1'b0}),
    .fci(\picorv32_core/add2/c31 ),
    .f({open_n20627,\picorv32_core/n450 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add2/ucin_al_u2538"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add2/u3_al_u2539  (
    .a({\picorv32_core/reg_pc [5],\picorv32_core/reg_pc [3]}),
    .b({\picorv32_core/reg_pc [6],\picorv32_core/reg_pc [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add2/c3 ),
    .f({\picorv32_core/n450 [5],\picorv32_core/n450 [3]}),
    .fco(\picorv32_core/add2/c7 ),
    .fx({\picorv32_core/n450 [6],\picorv32_core/n450 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add2/ucin_al_u2538"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add2/u7_al_u2540  (
    .a({\picorv32_core/reg_pc [9],\picorv32_core/reg_pc [7]}),
    .b({\picorv32_core/reg_pc [10],\picorv32_core/reg_pc [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add2/c7 ),
    .f({\picorv32_core/n450 [9],\picorv32_core/n450 [7]}),
    .fco(\picorv32_core/add2/c11 ),
    .fx({\picorv32_core/n450 [10],\picorv32_core/n450 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add2/ucin_al_u2538"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add2/ucin_al_u2538  (
    .a({\picorv32_core/reg_pc [1],1'b0}),
    .b({\picorv32_core/reg_pc [2],\picorv32_core/reg_pc [0]}),
    .c(2'b00),
    .d({\picorv32_core/latched_compr ,1'b1}),
    .e({\picorv32_core/n449 [2],1'b0}),
    .f({\picorv32_core/n450 [1],open_n20686}),
    .fco(\picorv32_core/add2/c3 ),
    .fx({\picorv32_core/n450 [2],\picorv32_core/n450 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u11_al_u2498  (
    .a({\picorv32_core/count_cycle [13],\picorv32_core/count_cycle [11]}),
    .b({\picorv32_core/count_cycle [14],\picorv32_core/count_cycle [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c11 ),
    .f({\picorv32_core/n459 [13],\picorv32_core/n459 [11]}),
    .fco(\picorv32_core/add3/c15 ),
    .fx({\picorv32_core/n459 [14],\picorv32_core/n459 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u15_al_u2499  (
    .a({\picorv32_core/count_cycle [17],\picorv32_core/count_cycle [15]}),
    .b({\picorv32_core/count_cycle [18],\picorv32_core/count_cycle [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c15 ),
    .f({\picorv32_core/n459 [17],\picorv32_core/n459 [15]}),
    .fco(\picorv32_core/add3/c19 ),
    .fx({\picorv32_core/n459 [18],\picorv32_core/n459 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u19_al_u2500  (
    .a({\picorv32_core/count_cycle [21],\picorv32_core/count_cycle [19]}),
    .b({\picorv32_core/count_cycle [22],\picorv32_core/count_cycle [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c19 ),
    .f({\picorv32_core/n459 [21],\picorv32_core/n459 [19]}),
    .fco(\picorv32_core/add3/c23 ),
    .fx({\picorv32_core/n459 [22],\picorv32_core/n459 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u23_al_u2501  (
    .a({\picorv32_core/count_cycle [25],\picorv32_core/count_cycle [23]}),
    .b({\picorv32_core/count_cycle [26],\picorv32_core/count_cycle [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c23 ),
    .f({\picorv32_core/n459 [25],\picorv32_core/n459 [23]}),
    .fco(\picorv32_core/add3/c27 ),
    .fx({\picorv32_core/n459 [26],\picorv32_core/n459 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u27_al_u2502  (
    .a({\picorv32_core/count_cycle [29],\picorv32_core/count_cycle [27]}),
    .b({\picorv32_core/count_cycle [30],\picorv32_core/count_cycle [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c27 ),
    .f({\picorv32_core/n459 [29],\picorv32_core/n459 [27]}),
    .fco(\picorv32_core/add3/c31 ),
    .fx({\picorv32_core/n459 [30],\picorv32_core/n459 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u31_al_u2503  (
    .a({\picorv32_core/count_cycle [33],\picorv32_core/count_cycle [31]}),
    .b({\picorv32_core/count_cycle [34],\picorv32_core/count_cycle [32]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c31 ),
    .f({\picorv32_core/n459 [33],\picorv32_core/n459 [31]}),
    .fco(\picorv32_core/add3/c35 ),
    .fx({\picorv32_core/n459 [34],\picorv32_core/n459 [32]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u35_al_u2504  (
    .a({\picorv32_core/count_cycle [37],\picorv32_core/count_cycle [35]}),
    .b({\picorv32_core/count_cycle [38],\picorv32_core/count_cycle [36]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c35 ),
    .f({\picorv32_core/n459 [37],\picorv32_core/n459 [35]}),
    .fco(\picorv32_core/add3/c39 ),
    .fx({\picorv32_core/n459 [38],\picorv32_core/n459 [36]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u39_al_u2505  (
    .a({\picorv32_core/count_cycle [41],\picorv32_core/count_cycle [39]}),
    .b({\picorv32_core/count_cycle [42],\picorv32_core/count_cycle [40]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c39 ),
    .f({\picorv32_core/n459 [41],\picorv32_core/n459 [39]}),
    .fco(\picorv32_core/add3/c43 ),
    .fx({\picorv32_core/n459 [42],\picorv32_core/n459 [40]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u3_al_u2496  (
    .a({\picorv32_core/count_cycle [5],\picorv32_core/count_cycle [3]}),
    .b({\picorv32_core/count_cycle [6],\picorv32_core/count_cycle [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c3 ),
    .f({\picorv32_core/n459 [5],\picorv32_core/n459 [3]}),
    .fco(\picorv32_core/add3/c7 ),
    .fx({\picorv32_core/n459 [6],\picorv32_core/n459 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u43_al_u2506  (
    .a({\picorv32_core/count_cycle [45],\picorv32_core/count_cycle [43]}),
    .b({\picorv32_core/count_cycle [46],\picorv32_core/count_cycle [44]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c43 ),
    .f({\picorv32_core/n459 [45],\picorv32_core/n459 [43]}),
    .fco(\picorv32_core/add3/c47 ),
    .fx({\picorv32_core/n459 [46],\picorv32_core/n459 [44]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y6Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u47_al_u2507  (
    .a({\picorv32_core/count_cycle [49],\picorv32_core/count_cycle [47]}),
    .b({\picorv32_core/count_cycle [50],\picorv32_core/count_cycle [48]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c47 ),
    .f({\picorv32_core/n459 [49],\picorv32_core/n459 [47]}),
    .fco(\picorv32_core/add3/c51 ),
    .fx({\picorv32_core/n459 [50],\picorv32_core/n459 [48]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y6Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u51_al_u2508  (
    .a({\picorv32_core/count_cycle [53],\picorv32_core/count_cycle [51]}),
    .b({\picorv32_core/count_cycle [54],\picorv32_core/count_cycle [52]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c51 ),
    .f({\picorv32_core/n459 [53],\picorv32_core/n459 [51]}),
    .fco(\picorv32_core/add3/c55 ),
    .fx({\picorv32_core/n459 [54],\picorv32_core/n459 [52]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y7Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u55_al_u2509  (
    .a({\picorv32_core/count_cycle [57],\picorv32_core/count_cycle [55]}),
    .b({\picorv32_core/count_cycle [58],\picorv32_core/count_cycle [56]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c55 ),
    .f({\picorv32_core/n459 [57],\picorv32_core/n459 [55]}),
    .fco(\picorv32_core/add3/c59 ),
    .fx({\picorv32_core/n459 [58],\picorv32_core/n459 [56]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y7Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u59_al_u2510  (
    .a({\picorv32_core/count_cycle [61],\picorv32_core/count_cycle [59]}),
    .b({\picorv32_core/count_cycle [62],\picorv32_core/count_cycle [60]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c59 ),
    .f({\picorv32_core/n459 [61],\picorv32_core/n459 [59]}),
    .fco(\picorv32_core/add3/c63 ),
    .fx({\picorv32_core/n459 [62],\picorv32_core/n459 [60]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y8Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u63_al_u2511  (
    .a({open_n20941,\picorv32_core/count_cycle [63]}),
    .c(2'b00),
    .d({open_n20946,1'b0}),
    .fci(\picorv32_core/add3/c63 ),
    .f({open_n20963,\picorv32_core/n459 [63]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add3/u7_al_u2497  (
    .a({\picorv32_core/count_cycle [9],\picorv32_core/count_cycle [7]}),
    .b({\picorv32_core/count_cycle [10],\picorv32_core/count_cycle [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add3/c7 ),
    .f({\picorv32_core/n459 [9],\picorv32_core/n459 [7]}),
    .fco(\picorv32_core/add3/c11 ),
    .fx({\picorv32_core/n459 [10],\picorv32_core/n459 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add3/ucin_al_u2495"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/add3/ucin_al_u2495  (
    .a({\picorv32_core/count_cycle [1],1'b0}),
    .b({\picorv32_core/count_cycle [2],\picorv32_core/count_cycle [0]}),
    .c(2'b00),
    .clk(clk_pad),
    .d(2'b01),
    .e(2'b01),
    .mi(\picorv32_core/n459 [1:0]),
    .sr(resetn_placeOpt_5),
    .f({\picorv32_core/n459 [1],open_n21000}),
    .fco(\picorv32_core/add3/c3 ),
    .fx({\picorv32_core/n459 [2],\picorv32_core/n459 [0]}),
    .q(\picorv32_core/count_cycle [1:0]));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add4/ucin_al_u2547"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add4/u11_al_u2550  (
    .a({\picorv32_core/n500 [13],\picorv32_core/n500 [11]}),
    .b({\picorv32_core/n500 [14],\picorv32_core/n500 [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add4/c11 ),
    .f({\picorv32_core/n502 [13],\picorv32_core/n502 [11]}),
    .fco(\picorv32_core/add4/c15 ),
    .fx({\picorv32_core/n502 [14],\picorv32_core/n502 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add4/ucin_al_u2547"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add4/u15_al_u2551  (
    .a({\picorv32_core/n500 [17],\picorv32_core/n500 [15]}),
    .b({\picorv32_core/n500 [18],\picorv32_core/n500 [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add4/c15 ),
    .f({\picorv32_core/n502 [17],\picorv32_core/n502 [15]}),
    .fco(\picorv32_core/add4/c19 ),
    .fx({\picorv32_core/n502 [18],\picorv32_core/n502 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add4/ucin_al_u2547"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add4/u19_al_u2552  (
    .a({\picorv32_core/n500 [21],\picorv32_core/n500 [19]}),
    .b({\picorv32_core/n500 [22],\picorv32_core/n500 [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add4/c19 ),
    .f({\picorv32_core/n502 [21],\picorv32_core/n502 [19]}),
    .fco(\picorv32_core/add4/c23 ),
    .fx({\picorv32_core/n502 [22],\picorv32_core/n502 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add4/ucin_al_u2547"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add4/u23_al_u2553  (
    .a({\picorv32_core/n500 [25],\picorv32_core/n500 [23]}),
    .b({\picorv32_core/n500 [26],\picorv32_core/n500 [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add4/c23 ),
    .f({\picorv32_core/n502 [25],\picorv32_core/n502 [23]}),
    .fco(\picorv32_core/add4/c27 ),
    .fx({\picorv32_core/n502 [26],\picorv32_core/n502 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add4/ucin_al_u2547"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add4/u27_al_u2554  (
    .a({\picorv32_core/n500 [29],\picorv32_core/n500 [27]}),
    .b({\picorv32_core/n500 [30],\picorv32_core/n500 [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add4/c27 ),
    .f({\picorv32_core/n502 [29],\picorv32_core/n502 [27]}),
    .fco(\picorv32_core/add4/c31 ),
    .fx({\picorv32_core/n502 [30],\picorv32_core/n502 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add4/ucin_al_u2547"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add4/u31_al_u2555  (
    .a({open_n21091,\picorv32_core/n500 [31]}),
    .c(2'b00),
    .d({open_n21096,1'b0}),
    .fci(\picorv32_core/add4/c31 ),
    .f({open_n21113,\picorv32_core/n502 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add4/ucin_al_u2547"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add4/u3_al_u2548  (
    .a({\picorv32_core/n500 [5],\picorv32_core/n500 [3]}),
    .b({\picorv32_core/n500 [6],\picorv32_core/n500 [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add4/c3 ),
    .f({\picorv32_core/n502 [5],\picorv32_core/n502 [3]}),
    .fco(\picorv32_core/add4/c7 ),
    .fx({\picorv32_core/n502 [6],\picorv32_core/n502 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add4/ucin_al_u2547"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add4/u7_al_u2549  (
    .a({\picorv32_core/n500 [9],\picorv32_core/n500 [7]}),
    .b({\picorv32_core/n500 [10],\picorv32_core/n500 [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add4/c7 ),
    .f({\picorv32_core/n502 [9],\picorv32_core/n502 [7]}),
    .fco(\picorv32_core/add4/c11 ),
    .fx({\picorv32_core/n502 [10],\picorv32_core/n502 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add4/ucin_al_u2547"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add4/ucin_al_u2547  (
    .a({\picorv32_core/n500 [1],1'b0}),
    .b({\picorv32_core/n500 [2],\picorv32_core/n500 [0]}),
    .c(2'b00),
    .d({\picorv32_core/compressed_instr ,1'b1}),
    .e({\picorv32_core/n501 [2],1'b0}),
    .f({\picorv32_core/n502 [1],open_n21172}),
    .fco(\picorv32_core/add4/c3 ),
    .fx({\picorv32_core/n502 [2],\picorv32_core/n502 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u11_al_u2515  (
    .a({\picorv32_core/count_instr [13],\picorv32_core/count_instr [11]}),
    .b({\picorv32_core/count_instr [14],\picorv32_core/count_instr [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c11 ),
    .f({\picorv32_core/n503 [13],\picorv32_core/n503 [11]}),
    .fco(\picorv32_core/add5/c15 ),
    .fx({\picorv32_core/n503 [14],\picorv32_core/n503 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u15_al_u2516  (
    .a({\picorv32_core/count_instr [17],\picorv32_core/count_instr [15]}),
    .b({\picorv32_core/count_instr [18],\picorv32_core/count_instr [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c15 ),
    .f({\picorv32_core/n503 [17],\picorv32_core/n503 [15]}),
    .fco(\picorv32_core/add5/c19 ),
    .fx({\picorv32_core/n503 [18],\picorv32_core/n503 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u19_al_u2517  (
    .a({\picorv32_core/count_instr [21],\picorv32_core/count_instr [19]}),
    .b({\picorv32_core/count_instr [22],\picorv32_core/count_instr [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c19 ),
    .f({\picorv32_core/n503 [21],\picorv32_core/n503 [19]}),
    .fco(\picorv32_core/add5/c23 ),
    .fx({\picorv32_core/n503 [22],\picorv32_core/n503 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u23_al_u2518  (
    .a({\picorv32_core/count_instr [25],\picorv32_core/count_instr [23]}),
    .b({\picorv32_core/count_instr [26],\picorv32_core/count_instr [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c23 ),
    .f({\picorv32_core/n503 [25],\picorv32_core/n503 [23]}),
    .fco(\picorv32_core/add5/c27 ),
    .fx({\picorv32_core/n503 [26],\picorv32_core/n503 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u27_al_u2519  (
    .a({\picorv32_core/count_instr [29],\picorv32_core/count_instr [27]}),
    .b({\picorv32_core/count_instr [30],\picorv32_core/count_instr [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c27 ),
    .f({\picorv32_core/n503 [29],\picorv32_core/n503 [27]}),
    .fco(\picorv32_core/add5/c31 ),
    .fx({\picorv32_core/n503 [30],\picorv32_core/n503 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u31_al_u2520  (
    .a({\picorv32_core/count_instr [33],\picorv32_core/count_instr [31]}),
    .b({\picorv32_core/count_instr [34],\picorv32_core/count_instr [32]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c31 ),
    .f({\picorv32_core/n503 [33],\picorv32_core/n503 [31]}),
    .fco(\picorv32_core/add5/c35 ),
    .fx({\picorv32_core/n503 [34],\picorv32_core/n503 [32]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u35_al_u2521  (
    .a({\picorv32_core/count_instr [37],\picorv32_core/count_instr [35]}),
    .b({\picorv32_core/count_instr [38],\picorv32_core/count_instr [36]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c35 ),
    .f({\picorv32_core/n503 [37],\picorv32_core/n503 [35]}),
    .fco(\picorv32_core/add5/c39 ),
    .fx({\picorv32_core/n503 [38],\picorv32_core/n503 [36]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u39_al_u2522  (
    .a({\picorv32_core/count_instr [41],\picorv32_core/count_instr [39]}),
    .b({\picorv32_core/count_instr [42],\picorv32_core/count_instr [40]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c39 ),
    .f({\picorv32_core/n503 [41],\picorv32_core/n503 [39]}),
    .fco(\picorv32_core/add5/c43 ),
    .fx({\picorv32_core/n503 [42],\picorv32_core/n503 [40]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u3_al_u2513  (
    .a({\picorv32_core/count_instr [5],\picorv32_core/count_instr [3]}),
    .b({\picorv32_core/count_instr [6],\picorv32_core/count_instr [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c3 ),
    .f({\picorv32_core/n503 [5],\picorv32_core/n503 [3]}),
    .fco(\picorv32_core/add5/c7 ),
    .fx({\picorv32_core/n503 [6],\picorv32_core/n503 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u43_al_u2523  (
    .a({\picorv32_core/count_instr [45],\picorv32_core/count_instr [43]}),
    .b({\picorv32_core/count_instr [46],\picorv32_core/count_instr [44]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c43 ),
    .f({\picorv32_core/n503 [45],\picorv32_core/n503 [43]}),
    .fco(\picorv32_core/add5/c47 ),
    .fx({\picorv32_core/n503 [46],\picorv32_core/n503 [44]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y6Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u47_al_u2524  (
    .a({\picorv32_core/count_instr [49],\picorv32_core/count_instr [47]}),
    .b({\picorv32_core/count_instr [50],\picorv32_core/count_instr [48]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c47 ),
    .f({\picorv32_core/n503 [49],\picorv32_core/n503 [47]}),
    .fco(\picorv32_core/add5/c51 ),
    .fx({\picorv32_core/n503 [50],\picorv32_core/n503 [48]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y6Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u51_al_u2525  (
    .a({\picorv32_core/count_instr [53],\picorv32_core/count_instr [51]}),
    .b({\picorv32_core/count_instr [54],\picorv32_core/count_instr [52]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c51 ),
    .f({\picorv32_core/n503 [53],\picorv32_core/n503 [51]}),
    .fco(\picorv32_core/add5/c55 ),
    .fx({\picorv32_core/n503 [54],\picorv32_core/n503 [52]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y7Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u55_al_u2526  (
    .a({\picorv32_core/count_instr [57],\picorv32_core/count_instr [55]}),
    .b({\picorv32_core/count_instr [58],\picorv32_core/count_instr [56]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c55 ),
    .f({\picorv32_core/n503 [57],\picorv32_core/n503 [55]}),
    .fco(\picorv32_core/add5/c59 ),
    .fx({\picorv32_core/n503 [58],\picorv32_core/n503 [56]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y7Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u59_al_u2527  (
    .a({\picorv32_core/count_instr [61],\picorv32_core/count_instr [59]}),
    .b({\picorv32_core/count_instr [62],\picorv32_core/count_instr [60]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c59 ),
    .f({\picorv32_core/n503 [61],\picorv32_core/n503 [59]}),
    .fco(\picorv32_core/add5/c63 ),
    .fx({\picorv32_core/n503 [62],\picorv32_core/n503 [60]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y8Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u63_al_u2528  (
    .a({open_n21427,\picorv32_core/count_instr [63]}),
    .c(2'b00),
    .d({open_n21432,1'b0}),
    .fci(\picorv32_core/add5/c63 ),
    .f({open_n21449,\picorv32_core/n503 [63]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add5/u7_al_u2514  (
    .a({\picorv32_core/count_instr [9],\picorv32_core/count_instr [7]}),
    .b({\picorv32_core/count_instr [10],\picorv32_core/count_instr [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\picorv32_core/add5/c7 ),
    .f({\picorv32_core/n503 [9],\picorv32_core/n503 [7]}),
    .fco(\picorv32_core/add5/c11 ),
    .fx({\picorv32_core/n503 [10],\picorv32_core/n503 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add5/ucin_al_u2512"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/add5/ucin_al_u2512  (
    .a({\picorv32_core/count_instr [1],1'b0}),
    .b({\picorv32_core/count_instr [2],\picorv32_core/count_instr [0]}),
    .c(2'b00),
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d(2'b01),
    .e(2'b01),
    .mi(\picorv32_core/n503 [1:0]),
    .sr(resetn_placeOpt_5),
    .f({\picorv32_core/n503 [1],open_n21485}),
    .fco(\picorv32_core/add5/c3 ),
    .fx({\picorv32_core/n503 [2],\picorv32_core/n503 [0]}),
    .q(\picorv32_core/count_instr [1:0]));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add6/ucin_al_u2556"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add6/u11_al_u2559  (
    .a({\picorv32_core/n500 [13],\picorv32_core/n500 [11]}),
    .b({\picorv32_core/n500 [14],\picorv32_core/n500 [12]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm_uj [13],\picorv32_core/decoded_imm_uj [11]}),
    .e({\picorv32_core/decoded_imm_uj [14],\picorv32_core/decoded_imm_uj [12]}),
    .fci(\picorv32_core/add6/c11 ),
    .f({\picorv32_core/n504 [13],\picorv32_core/n504 [11]}),
    .fco(\picorv32_core/add6/c15 ),
    .fx({\picorv32_core/n504 [14],\picorv32_core/n504 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add6/ucin_al_u2556"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add6/u15_al_u2560  (
    .a({\picorv32_core/n500 [17],\picorv32_core/n500 [15]}),
    .b({\picorv32_core/n500 [18],\picorv32_core/n500 [16]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm_uj [17],\picorv32_core/decoded_imm_uj [15]}),
    .e({\picorv32_core/decoded_imm_uj [18],\picorv32_core/decoded_imm_uj [16]}),
    .fci(\picorv32_core/add6/c15 ),
    .f({\picorv32_core/n504 [17],\picorv32_core/n504 [15]}),
    .fco(\picorv32_core/add6/c19 ),
    .fx({\picorv32_core/n504 [18],\picorv32_core/n504 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add6/ucin_al_u2556"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add6/u19_al_u2561  (
    .a({\picorv32_core/n500 [21],\picorv32_core/n500 [19]}),
    .b({\picorv32_core/n500 [22],\picorv32_core/n500 [20]}),
    .c(2'b00),
    .d(\picorv32_core/decoded_imm_uj [20:19]),
    .e({\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20]}),
    .fci(\picorv32_core/add6/c19 ),
    .f({\picorv32_core/n504 [21],\picorv32_core/n504 [19]}),
    .fco(\picorv32_core/add6/c23 ),
    .fx({\picorv32_core/n504 [22],\picorv32_core/n504 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add6/ucin_al_u2556"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add6/u23_al_u2562  (
    .a({\picorv32_core/n500 [25],\picorv32_core/n500 [23]}),
    .b({\picorv32_core/n500 [26],\picorv32_core/n500 [24]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20]}),
    .e({\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20]}),
    .fci(\picorv32_core/add6/c23 ),
    .f({\picorv32_core/n504 [25],\picorv32_core/n504 [23]}),
    .fco(\picorv32_core/add6/c27 ),
    .fx({\picorv32_core/n504 [26],\picorv32_core/n504 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add6/ucin_al_u2556"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add6/u27_al_u2563  (
    .a({\picorv32_core/n500 [29],\picorv32_core/n500 [27]}),
    .b({\picorv32_core/n500 [30],\picorv32_core/n500 [28]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20]}),
    .e({\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20]}),
    .fci(\picorv32_core/add6/c27 ),
    .f({\picorv32_core/n504 [29],\picorv32_core/n504 [27]}),
    .fco(\picorv32_core/add6/c31 ),
    .fx({\picorv32_core/n504 [30],\picorv32_core/n504 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add6/ucin_al_u2556"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add6/u31_al_u2564  (
    .a({open_n21576,\picorv32_core/n500 [31]}),
    .c(2'b00),
    .d({open_n21581,\picorv32_core/decoded_imm_uj [20]}),
    .fci(\picorv32_core/add6/c31 ),
    .f({open_n21598,\picorv32_core/n504 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add6/ucin_al_u2556"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add6/u3_al_u2557  (
    .a({\picorv32_core/n500 [5],\picorv32_core/n500 [3]}),
    .b({\picorv32_core/n500 [6],\picorv32_core/n500 [4]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm_uj [5],\picorv32_core/decoded_imm_uj [3]}),
    .e({\picorv32_core/decoded_imm_uj [6],\picorv32_core/decoded_imm_uj [4]}),
    .fci(\picorv32_core/add6/c3 ),
    .f({\picorv32_core/n504 [5],\picorv32_core/n504 [3]}),
    .fco(\picorv32_core/add6/c7 ),
    .fx({\picorv32_core/n504 [6],\picorv32_core/n504 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add6/ucin_al_u2556"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add6/u7_al_u2558  (
    .a({\picorv32_core/n500 [9],\picorv32_core/n500 [7]}),
    .b({\picorv32_core/n500 [10],\picorv32_core/n500 [8]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm_uj [9],\picorv32_core/decoded_imm_uj [7]}),
    .e({\picorv32_core/decoded_imm_uj [10],\picorv32_core/decoded_imm_uj [8]}),
    .fci(\picorv32_core/add6/c7 ),
    .f({\picorv32_core/n504 [9],\picorv32_core/n504 [7]}),
    .fco(\picorv32_core/add6/c11 ),
    .fx({\picorv32_core/n504 [10],\picorv32_core/n504 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add6/ucin_al_u2556"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add6/ucin_al_u2556  (
    .a({\picorv32_core/n500 [1],1'b0}),
    .b({\picorv32_core/n500 [2],\picorv32_core/n500 [0]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm_uj [1],1'b1}),
    .e({\picorv32_core/decoded_imm_uj [2],1'b0}),
    .f({\picorv32_core/n504 [1],open_n21657}),
    .fco(\picorv32_core/add6/c3 ),
    .fx({\picorv32_core/n504 [2],\picorv32_core/n504 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add7/ucin_al_u2565"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add7/u11_al_u2568  (
    .a({\picorv32_core/reg_pc [13],\picorv32_core/reg_pc [11]}),
    .b({\picorv32_core/reg_pc [14],\picorv32_core/reg_pc [12]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm [13],\picorv32_core/decoded_imm [11]}),
    .e({\picorv32_core/decoded_imm [14],\picorv32_core/decoded_imm [12]}),
    .fci(\picorv32_core/add7/c11 ),
    .f({\picorv32_core/n543 [13],\picorv32_core/n543 [11]}),
    .fco(\picorv32_core/add7/c15 ),
    .fx({\picorv32_core/n543 [14],\picorv32_core/n543 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add7/ucin_al_u2565"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add7/u15_al_u2569  (
    .a({\picorv32_core/reg_pc [17],\picorv32_core/reg_pc [15]}),
    .b({\picorv32_core/reg_pc [18],\picorv32_core/reg_pc [16]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm [17],\picorv32_core/decoded_imm [15]}),
    .e({\picorv32_core/decoded_imm [18],\picorv32_core/decoded_imm [16]}),
    .fci(\picorv32_core/add7/c15 ),
    .f({\picorv32_core/n543 [17],\picorv32_core/n543 [15]}),
    .fco(\picorv32_core/add7/c19 ),
    .fx({\picorv32_core/n543 [18],\picorv32_core/n543 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add7/ucin_al_u2565"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add7/u19_al_u2570  (
    .a({\picorv32_core/reg_pc [21],\picorv32_core/reg_pc [19]}),
    .b({\picorv32_core/reg_pc [22],\picorv32_core/reg_pc [20]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm [21],\picorv32_core/decoded_imm [19]}),
    .e({\picorv32_core/decoded_imm [22],\picorv32_core/decoded_imm [20]}),
    .fci(\picorv32_core/add7/c19 ),
    .f({\picorv32_core/n543 [21],\picorv32_core/n543 [19]}),
    .fco(\picorv32_core/add7/c23 ),
    .fx({\picorv32_core/n543 [22],\picorv32_core/n543 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add7/ucin_al_u2565"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add7/u23_al_u2571  (
    .a({\picorv32_core/reg_pc [25],\picorv32_core/reg_pc [23]}),
    .b({\picorv32_core/reg_pc [26],\picorv32_core/reg_pc [24]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm [25],\picorv32_core/decoded_imm [23]}),
    .e({\picorv32_core/decoded_imm [26],\picorv32_core/decoded_imm [24]}),
    .fci(\picorv32_core/add7/c23 ),
    .f({\picorv32_core/n543 [25],\picorv32_core/n543 [23]}),
    .fco(\picorv32_core/add7/c27 ),
    .fx({\picorv32_core/n543 [26],\picorv32_core/n543 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add7/ucin_al_u2565"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add7/u27_al_u2572  (
    .a({\picorv32_core/reg_pc [29],\picorv32_core/reg_pc [27]}),
    .b({\picorv32_core/reg_pc [30],\picorv32_core/reg_pc [28]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm [29],\picorv32_core/decoded_imm [27]}),
    .e({\picorv32_core/decoded_imm [30],\picorv32_core/decoded_imm [28]}),
    .fci(\picorv32_core/add7/c27 ),
    .f({\picorv32_core/n543 [29],\picorv32_core/n543 [27]}),
    .fco(\picorv32_core/add7/c31 ),
    .fx({\picorv32_core/n543 [30],\picorv32_core/n543 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add7/ucin_al_u2565"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add7/u31_al_u2573  (
    .a({open_n21750,\picorv32_core/reg_pc [31]}),
    .c(2'b00),
    .d({open_n21755,\picorv32_core/decoded_imm [31]}),
    .fci(\picorv32_core/add7/c31 ),
    .f({open_n21772,\picorv32_core/n543 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add7/ucin_al_u2565"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add7/u3_al_u2566  (
    .a({\picorv32_core/reg_pc [5],\picorv32_core/reg_pc [3]}),
    .b({\picorv32_core/reg_pc [6],\picorv32_core/reg_pc [4]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm [5],\picorv32_core/decoded_imm [3]}),
    .e({\picorv32_core/decoded_imm [6],\picorv32_core/decoded_imm [4]}),
    .fci(\picorv32_core/add7/c3 ),
    .f({\picorv32_core/n543 [5],\picorv32_core/n543 [3]}),
    .fco(\picorv32_core/add7/c7 ),
    .fx({\picorv32_core/n543 [6],\picorv32_core/n543 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add7/ucin_al_u2565"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add7/u7_al_u2567  (
    .a({\picorv32_core/reg_pc [9],\picorv32_core/reg_pc [7]}),
    .b({\picorv32_core/reg_pc [10],\picorv32_core/reg_pc [8]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm [9],\picorv32_core/decoded_imm [7]}),
    .e({\picorv32_core/decoded_imm [10],\picorv32_core/decoded_imm [8]}),
    .fci(\picorv32_core/add7/c7 ),
    .f({\picorv32_core/n543 [9],\picorv32_core/n543 [7]}),
    .fco(\picorv32_core/add7/c11 ),
    .fx({\picorv32_core/n543 [10],\picorv32_core/n543 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/add7/ucin_al_u2565"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \picorv32_core/add7/ucin_al_u2565  (
    .a({\picorv32_core/reg_pc [1],1'b0}),
    .b({\picorv32_core/reg_pc [2],\picorv32_core/reg_pc [0]}),
    .c(2'b00),
    .d({\picorv32_core/decoded_imm [1],1'b1}),
    .e({\picorv32_core/decoded_imm [2],\picorv32_core/decoded_imm [0]}),
    .f({\picorv32_core/n543 [1],open_n21831}),
    .fco(\picorv32_core/add7/c3 ),
    .fx({\picorv32_core/n543 [2],\picorv32_core/n543 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u0|picorv32_core/add8/ucin  (
    .a({\picorv32_core/pcpi_rs1$0$ ,1'b0}),
    .b({\picorv32_core/decoded_imm [0],open_n21834}),
    .f({\picorv32_core/n576 [0],open_n21854}),
    .fco(\picorv32_core/add8/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u10|picorv32_core/add8/u9  (
    .a({\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$9$ }),
    .b(\picorv32_core/decoded_imm [10:9]),
    .fci(\picorv32_core/add8/c9 ),
    .f(\picorv32_core/n576 [10:9]),
    .fco(\picorv32_core/add8/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u12|picorv32_core/add8/u11  (
    .a({\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/pcpi_rs1$11$ }),
    .b(\picorv32_core/decoded_imm [12:11]),
    .fci(\picorv32_core/add8/c11 ),
    .f(\picorv32_core/n576 [12:11]),
    .fco(\picorv32_core/add8/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u14|picorv32_core/add8/u13  (
    .a({\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$13$ }),
    .b(\picorv32_core/decoded_imm [14:13]),
    .fci(\picorv32_core/add8/c13 ),
    .f(\picorv32_core/n576 [14:13]),
    .fco(\picorv32_core/add8/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u16|picorv32_core/add8/u15  (
    .a({\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/pcpi_rs1$15$ }),
    .b(\picorv32_core/decoded_imm [16:15]),
    .fci(\picorv32_core/add8/c15 ),
    .f(\picorv32_core/n576 [16:15]),
    .fco(\picorv32_core/add8/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u18|picorv32_core/add8/u17  (
    .a({\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$17$ }),
    .b(\picorv32_core/decoded_imm [18:17]),
    .fci(\picorv32_core/add8/c17 ),
    .f(\picorv32_core/n576 [18:17]),
    .fco(\picorv32_core/add8/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u20|picorv32_core/add8/u19  (
    .a({\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/pcpi_rs1$19$ }),
    .b(\picorv32_core/decoded_imm [20:19]),
    .fci(\picorv32_core/add8/c19 ),
    .f(\picorv32_core/n576 [20:19]),
    .fco(\picorv32_core/add8/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u22|picorv32_core/add8/u21  (
    .a({\picorv32_core/decoded_imm [22],\picorv32_core/pcpi_rs1$21$ }),
    .b({\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/decoded_imm [21]}),
    .fci(\picorv32_core/add8/c21 ),
    .f(\picorv32_core/n576 [22:21]),
    .fco(\picorv32_core/add8/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u24|picorv32_core/add8/u23  (
    .a({\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/pcpi_rs1$23$ }),
    .b(\picorv32_core/decoded_imm [24:23]),
    .fci(\picorv32_core/add8/c23 ),
    .f(\picorv32_core/n576 [24:23]),
    .fco(\picorv32_core/add8/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u26|picorv32_core/add8/u25  (
    .a({\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$25$ }),
    .b(\picorv32_core/decoded_imm [26:25]),
    .fci(\picorv32_core/add8/c25 ),
    .f(\picorv32_core/n576 [26:25]),
    .fco(\picorv32_core/add8/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u28|picorv32_core/add8/u27  (
    .a({\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/pcpi_rs1$27$ }),
    .b(\picorv32_core/decoded_imm [28:27]),
    .fci(\picorv32_core/add8/c27 ),
    .f(\picorv32_core/n576 [28:27]),
    .fco(\picorv32_core/add8/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u2|picorv32_core/add8/u1  (
    .a({\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$1$ }),
    .b(\picorv32_core/decoded_imm [2:1]),
    .fci(\picorv32_core/add8/c1 ),
    .f(\picorv32_core/n576 [2:1]),
    .fco(\picorv32_core/add8/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u30|picorv32_core/add8/u29  (
    .a({\picorv32_core/pcpi_rs1$30$ ,\picorv32_core/pcpi_rs1$29$ }),
    .b(\picorv32_core/decoded_imm [30:29]),
    .fci(\picorv32_core/add8/c29 ),
    .f(\picorv32_core/n576 [30:29]),
    .fco(\picorv32_core/add8/c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u31_al_u2575  (
    .a({open_n22123,\picorv32_core/pcpi_rs1$31$ }),
    .b({open_n22124,\picorv32_core/decoded_imm [31]}),
    .fci(\picorv32_core/add8/c31 ),
    .f({open_n22143,\picorv32_core/n576 [31]}));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u4|picorv32_core/add8/u3  (
    .a({\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/pcpi_rs1$3$ }),
    .b(\picorv32_core/decoded_imm [4:3]),
    .fci(\picorv32_core/add8/c3 ),
    .f(\picorv32_core/n576 [4:3]),
    .fco(\picorv32_core/add8/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u6|picorv32_core/add8/u5  (
    .a({\picorv32_core/pcpi_rs1$6$ ,\picorv32_core/pcpi_rs1$5$ }),
    .b(\picorv32_core/decoded_imm [6:5]),
    .fci(\picorv32_core/add8/c5 ),
    .f(\picorv32_core/n576 [6:5]),
    .fco(\picorv32_core/add8/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/add8/u0|picorv32_core/add8/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \picorv32_core/add8/u8|picorv32_core/add8/u7  (
    .a({\picorv32_core/decoded_imm [8],\picorv32_core/pcpi_rs1$7$ }),
    .b({\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/decoded_imm [7]}),
    .fci(\picorv32_core/add8/c7 ),
    .f(\picorv32_core/n576 [8:7]),
    .fco(\picorv32_core/add8/c9 ));
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*D*~(C*~(~0*B)))"),
    //.LUT1("~(~A*C*~(D*~(~1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101011111111),
    .INIT_LUT1(16'b1111111110101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/compressed_instr_reg  (
    .a({_al_u1296_o,_al_u1296_o}),
    .b({\picorv32_core/mem_rdata_latched_noshuffle [1],\picorv32_core/mem_rdata_latched_noshuffle [1]}),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_3 ,_al_u1295_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u1295_o,\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }),
    .mi({open_n22225,_al_u1088_o}),
    .fx({open_n22230,\picorv32_core/n180 }),
    .q({open_n22231,\picorv32_core/compressed_instr }));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c0_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r0_c0_l  (
    .a({\picorv32_core/cpuregs_wrdata [0],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [1],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [2],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [3],\picorv32_core/latched_rd [3]}),
    .e({open_n22233,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c0_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c0_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c0_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c0_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c0_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c0_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c0_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c0_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c0_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c0_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c0_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c0_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_001 ,\picorv32_core/cpuregs_p1/dram_do_i0_000 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c0_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c0_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c0_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c0_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c0_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c0_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c0_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_003 ,\picorv32_core/cpuregs_p1/dram_do_i0_002 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c1_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r0_c1_l  (
    .a({\picorv32_core/cpuregs_wrdata [4],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [5],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [6],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [7],\picorv32_core/latched_rd [3]}),
    .e({open_n22268,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c1_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c1_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c1_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c1_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c1_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c1_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c1_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c1_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c1_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c1_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c1_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c1_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_005 ,\picorv32_core/cpuregs_p1/dram_do_i0_004 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c1_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c1_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c1_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c1_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c1_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c1_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c1_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_007 ,\picorv32_core/cpuregs_p1/dram_do_i0_006 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c2_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r0_c2_l  (
    .a({\picorv32_core/cpuregs_wrdata [8],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [9],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [10],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [11],\picorv32_core/latched_rd [3]}),
    .e({open_n22303,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c2_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c2_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c2_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c2_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c2_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c2_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c2_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c2_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c2_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c2_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c2_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c2_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_009 ,\picorv32_core/cpuregs_p1/dram_do_i0_008 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c2_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c2_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c2_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c2_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c2_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c2_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c2_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_011 ,\picorv32_core/cpuregs_p1/dram_do_i0_010 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c3_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r0_c3_l  (
    .a({\picorv32_core/cpuregs_wrdata [12],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [13],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [14],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [15],\picorv32_core/latched_rd [3]}),
    .e({open_n22338,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c3_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c3_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c3_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c3_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c3_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c3_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c3_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c3_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c3_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c3_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c3_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c3_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_013 ,\picorv32_core/cpuregs_p1/dram_do_i0_012 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c3_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c3_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c3_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c3_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c3_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c3_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c3_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_015 ,\picorv32_core/cpuregs_p1/dram_do_i0_014 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c4_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r0_c4_l  (
    .a({\picorv32_core/cpuregs_wrdata [16],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [17],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [18],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [19],\picorv32_core/latched_rd [3]}),
    .e({open_n22373,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c4_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c4_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c4_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c4_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c4_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c4_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c4_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c4_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c4_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c4_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c4_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c4_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_017 ,\picorv32_core/cpuregs_p1/dram_do_i0_016 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c4_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c4_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c4_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c4_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c4_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c4_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c4_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_019 ,\picorv32_core/cpuregs_p1/dram_do_i0_018 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c5_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r0_c5_l  (
    .a({\picorv32_core/cpuregs_wrdata [20],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [21],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [22],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [23],\picorv32_core/latched_rd [3]}),
    .e({open_n22408,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c5_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c5_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c5_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c5_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c5_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c5_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c5_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c5_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c5_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c5_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c5_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c5_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_021 ,\picorv32_core/cpuregs_p1/dram_do_i0_020 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c5_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c5_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c5_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c5_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c5_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c5_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c5_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_023 ,\picorv32_core/cpuregs_p1/dram_do_i0_022 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c6_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r0_c6_l  (
    .a({\picorv32_core/cpuregs_wrdata [24],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [25],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [26],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [27],\picorv32_core/latched_rd [3]}),
    .e({open_n22443,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c6_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c6_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c6_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c6_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c6_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c6_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c6_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c6_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c6_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c6_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c6_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c6_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_025 ,\picorv32_core/cpuregs_p1/dram_do_i0_024 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c6_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c6_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c6_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c6_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c6_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c6_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c6_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_027 ,\picorv32_core/cpuregs_p1/dram_do_i0_026 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c7_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r0_c7_l  (
    .a({\picorv32_core/cpuregs_wrdata [28],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [29],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [30],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [31],\picorv32_core/latched_rd [3]}),
    .e({open_n22478,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c7_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c7_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c7_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c7_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c7_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c7_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c7_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c7_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c7_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c7_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c7_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c7_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_029 ,\picorv32_core/cpuregs_p1/dram_do_i0_028 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r0_c7_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r0_c7_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r0_c7_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r0_c7_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r0_c7_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r0_c7_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r0_c7_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i0_031 ,\picorv32_core/cpuregs_p1/dram_do_i0_030 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c0_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r1_c0_l  (
    .a({\picorv32_core/cpuregs_wrdata [0],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [1],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [2],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [3],\picorv32_core/latched_rd [3]}),
    .e({open_n22513,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c0_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c0_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c0_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c0_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c0_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c0_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c0_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c0_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c0_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c0_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c0_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c0_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_001 ,\picorv32_core/cpuregs_p1/dram_do_i1_000 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c0_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c0_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c0_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c0_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c0_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c0_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c0_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_003 ,\picorv32_core/cpuregs_p1/dram_do_i1_002 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c1_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r1_c1_l  (
    .a({\picorv32_core/cpuregs_wrdata [4],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [5],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [6],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [7],\picorv32_core/latched_rd [3]}),
    .e({open_n22548,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c1_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c1_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c1_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c1_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c1_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c1_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c1_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c1_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c1_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c1_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c1_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c1_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_005 ,\picorv32_core/cpuregs_p1/dram_do_i1_004 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c1_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c1_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c1_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c1_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c1_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c1_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c1_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_007 ,\picorv32_core/cpuregs_p1/dram_do_i1_006 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c2_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r1_c2_l  (
    .a({\picorv32_core/cpuregs_wrdata [8],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [9],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [10],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [11],\picorv32_core/latched_rd [3]}),
    .e({open_n22583,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c2_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c2_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c2_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c2_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c2_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c2_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c2_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c2_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c2_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c2_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c2_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c2_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_009 ,\picorv32_core/cpuregs_p1/dram_do_i1_008 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c2_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c2_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c2_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c2_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c2_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c2_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c2_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_011 ,\picorv32_core/cpuregs_p1/dram_do_i1_010 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c3_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r1_c3_l  (
    .a({\picorv32_core/cpuregs_wrdata [12],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [13],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [14],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [15],\picorv32_core/latched_rd [3]}),
    .e({open_n22618,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c3_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c3_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c3_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c3_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c3_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c3_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c3_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c3_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c3_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c3_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c3_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c3_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_013 ,\picorv32_core/cpuregs_p1/dram_do_i1_012 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c3_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c3_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c3_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c3_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c3_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c3_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c3_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_015 ,\picorv32_core/cpuregs_p1/dram_do_i1_014 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c4_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r1_c4_l  (
    .a({\picorv32_core/cpuregs_wrdata [16],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [17],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [18],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [19],\picorv32_core/latched_rd [3]}),
    .e({open_n22653,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c4_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c4_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c4_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c4_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c4_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c4_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c4_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c4_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c4_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c4_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c4_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c4_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_017 ,\picorv32_core/cpuregs_p1/dram_do_i1_016 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c4_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c4_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c4_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c4_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c4_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c4_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c4_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_019 ,\picorv32_core/cpuregs_p1/dram_do_i1_018 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c5_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r1_c5_l  (
    .a({\picorv32_core/cpuregs_wrdata [20],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [21],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [22],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [23],\picorv32_core/latched_rd [3]}),
    .e({open_n22688,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c5_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c5_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c5_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c5_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c5_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c5_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c5_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c5_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c5_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c5_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c5_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c5_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_021 ,\picorv32_core/cpuregs_p1/dram_do_i1_020 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c5_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c5_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c5_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c5_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c5_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c5_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c5_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_023 ,\picorv32_core/cpuregs_p1/dram_do_i1_022 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c6_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r1_c6_l  (
    .a({\picorv32_core/cpuregs_wrdata [24],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [25],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [26],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [27],\picorv32_core/latched_rd [3]}),
    .e({open_n22723,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c6_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c6_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c6_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c6_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c6_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c6_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c6_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c6_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c6_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c6_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c6_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c6_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_025 ,\picorv32_core/cpuregs_p1/dram_do_i1_024 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c6_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c6_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c6_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c6_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c6_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c6_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c6_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_027 ,\picorv32_core/cpuregs_p1/dram_do_i1_026 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c7_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p1/dram_r1_c7_l  (
    .a({\picorv32_core/cpuregs_wrdata [28],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [29],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [30],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [31],\picorv32_core/latched_rd [3]}),
    .e({open_n22758,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c7_di ),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c7_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c7_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c7_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c7_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c7_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c7_m0  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c7_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c7_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c7_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c7_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c7_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_029 ,\picorv32_core/cpuregs_p1/dram_do_i1_028 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p1/dram_r1_c7_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p1/dram_r1_c7_m1  (
    .a({\picorv32_core/decoded_rs1 [0],\picorv32_core/decoded_rs1 [0]}),
    .b({\picorv32_core/decoded_rs1 [1],\picorv32_core/decoded_rs1 [1]}),
    .c({\picorv32_core/decoded_rs1 [2],\picorv32_core/decoded_rs1 [2]}),
    .d({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_rs1 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p1/dram_r1_c7_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p1/dram_r1_c7_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p1/dram_r1_c7_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p1/dram_r1_c7_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p1/dram_r1_c7_we ),
    .f({\picorv32_core/cpuregs_p1/dram_do_i1_031 ,\picorv32_core/cpuregs_p1/dram_do_i1_030 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c0_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r0_c0_l  (
    .a({\picorv32_core/cpuregs_wrdata [0],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [1],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [2],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [3],\picorv32_core/latched_rd [3]}),
    .e({open_n22793,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c0_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c0_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c0_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c0_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c0_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c0_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c0_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c0_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c0_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c0_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c0_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c0_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_001 ,\picorv32_core/cpuregs_p2/dram_do_i0_000 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c0_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c0_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c0_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c0_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c0_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c0_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c0_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_003 ,\picorv32_core/cpuregs_p2/dram_do_i0_002 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c1_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r0_c1_l  (
    .a({\picorv32_core/cpuregs_wrdata [4],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [5],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [6],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [7],\picorv32_core/latched_rd [3]}),
    .e({open_n22828,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c1_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c1_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c1_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c1_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c1_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c1_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c1_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c1_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c1_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c1_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c1_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c1_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_005 ,\picorv32_core/cpuregs_p2/dram_do_i0_004 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c1_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c1_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c1_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c1_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c1_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c1_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c1_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_007 ,\picorv32_core/cpuregs_p2/dram_do_i0_006 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c2_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r0_c2_l  (
    .a({\picorv32_core/cpuregs_wrdata [8],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [9],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [10],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [11],\picorv32_core/latched_rd [3]}),
    .e({open_n22863,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c2_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c2_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c2_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c2_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c2_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c2_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c2_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c2_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c2_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c2_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c2_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c2_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_009 ,\picorv32_core/cpuregs_p2/dram_do_i0_008 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c2_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c2_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c2_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c2_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c2_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c2_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c2_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_011 ,\picorv32_core/cpuregs_p2/dram_do_i0_010 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c3_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r0_c3_l  (
    .a({\picorv32_core/cpuregs_wrdata [12],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [13],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [14],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [15],\picorv32_core/latched_rd [3]}),
    .e({open_n22898,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c3_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c3_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c3_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c3_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c3_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c3_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c3_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c3_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c3_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c3_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c3_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c3_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_013 ,\picorv32_core/cpuregs_p2/dram_do_i0_012 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c3_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c3_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c3_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c3_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c3_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c3_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c3_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_015 ,\picorv32_core/cpuregs_p2/dram_do_i0_014 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c4_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r0_c4_l  (
    .a({\picorv32_core/cpuregs_wrdata [16],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [17],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [18],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [19],\picorv32_core/latched_rd [3]}),
    .e({open_n22933,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c4_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c4_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c4_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c4_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c4_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c4_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c4_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c4_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c4_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c4_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c4_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c4_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_017 ,\picorv32_core/cpuregs_p2/dram_do_i0_016 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c4_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c4_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c4_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c4_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c4_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c4_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c4_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_019 ,\picorv32_core/cpuregs_p2/dram_do_i0_018 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c5_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r0_c5_l  (
    .a({\picorv32_core/cpuregs_wrdata [20],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [21],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [22],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [23],\picorv32_core/latched_rd [3]}),
    .e({open_n22968,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c5_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c5_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c5_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c5_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c5_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c5_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c5_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c5_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c5_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c5_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c5_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c5_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_021 ,\picorv32_core/cpuregs_p2/dram_do_i0_020 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c5_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c5_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c5_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c5_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c5_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c5_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c5_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_023 ,\picorv32_core/cpuregs_p2/dram_do_i0_022 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c6_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r0_c6_l  (
    .a({\picorv32_core/cpuregs_wrdata [24],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [25],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [26],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [27],\picorv32_core/latched_rd [3]}),
    .e({open_n23003,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c6_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c6_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c6_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c6_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c6_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c6_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c6_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c6_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c6_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c6_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c6_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c6_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_025 ,\picorv32_core/cpuregs_p2/dram_do_i0_024 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c6_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c6_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c6_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c6_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c6_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c6_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c6_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_027 ,\picorv32_core/cpuregs_p2/dram_do_i0_026 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c7_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r0_c7_l  (
    .a({\picorv32_core/cpuregs_wrdata [28],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [29],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [30],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [31],\picorv32_core/latched_rd [3]}),
    .e({open_n23038,\picorv32_core/n456_0_al_n603 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c7_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c7_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c7_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c7_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c7_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c7_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c7_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c7_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c7_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c7_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c7_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c7_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_029 ,\picorv32_core/cpuregs_p2/dram_do_i0_028 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r0_c7_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r0_c7_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r0_c7_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r0_c7_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r0_c7_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r0_c7_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r0_c7_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i0_031 ,\picorv32_core/cpuregs_p2/dram_do_i0_030 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c0_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r1_c0_l  (
    .a({\picorv32_core/cpuregs_wrdata [0],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [1],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [2],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [3],\picorv32_core/latched_rd [3]}),
    .e({open_n23073,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c0_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c0_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c0_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c0_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c0_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c0_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c0_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c0_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c0_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c0_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c0_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c0_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_001 ,\picorv32_core/cpuregs_p2/dram_do_i1_000 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c0_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c0_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c0_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c0_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c0_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c0_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c0_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_003 ,\picorv32_core/cpuregs_p2/dram_do_i1_002 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c1_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r1_c1_l  (
    .a({\picorv32_core/cpuregs_wrdata [4],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [5],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [6],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [7],\picorv32_core/latched_rd [3]}),
    .e({open_n23108,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c1_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c1_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c1_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c1_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c1_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c1_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c1_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c1_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c1_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c1_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c1_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c1_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_005 ,\picorv32_core/cpuregs_p2/dram_do_i1_004 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c1_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c1_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c1_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c1_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c1_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c1_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c1_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_007 ,\picorv32_core/cpuregs_p2/dram_do_i1_006 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c2_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r1_c2_l  (
    .a({\picorv32_core/cpuregs_wrdata [8],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [9],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [10],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [11],\picorv32_core/latched_rd [3]}),
    .e({open_n23143,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c2_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c2_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c2_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c2_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c2_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c2_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c2_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c2_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c2_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c2_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c2_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c2_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_009 ,\picorv32_core/cpuregs_p2/dram_do_i1_008 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c2_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c2_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c2_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c2_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c2_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c2_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c2_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_011 ,\picorv32_core/cpuregs_p2/dram_do_i1_010 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c3_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r1_c3_l  (
    .a({\picorv32_core/cpuregs_wrdata [12],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [13],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [14],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [15],\picorv32_core/latched_rd [3]}),
    .e({open_n23178,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c3_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c3_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c3_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c3_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c3_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c3_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c3_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c3_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c3_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c3_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c3_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c3_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_013 ,\picorv32_core/cpuregs_p2/dram_do_i1_012 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c3_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c3_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c3_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c3_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c3_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c3_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c3_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_015 ,\picorv32_core/cpuregs_p2/dram_do_i1_014 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c4_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r1_c4_l  (
    .a({\picorv32_core/cpuregs_wrdata [16],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [17],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [18],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [19],\picorv32_core/latched_rd [3]}),
    .e({open_n23213,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c4_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c4_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c4_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c4_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c4_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c4_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c4_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c4_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c4_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c4_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c4_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c4_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_017 ,\picorv32_core/cpuregs_p2/dram_do_i1_016 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c4_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c4_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c4_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c4_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c4_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c4_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c4_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_019 ,\picorv32_core/cpuregs_p2/dram_do_i1_018 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c5_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r1_c5_l  (
    .a({\picorv32_core/cpuregs_wrdata [20],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [21],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [22],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [23],\picorv32_core/latched_rd [3]}),
    .e({open_n23248,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c5_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c5_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c5_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c5_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c5_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c5_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c5_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c5_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c5_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c5_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c5_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c5_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_021 ,\picorv32_core/cpuregs_p2/dram_do_i1_020 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c5_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c5_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c5_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c5_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c5_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c5_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c5_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_023 ,\picorv32_core/cpuregs_p2/dram_do_i1_022 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c6_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r1_c6_l  (
    .a({\picorv32_core/cpuregs_wrdata [24],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [25],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [26],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [27],\picorv32_core/latched_rd [3]}),
    .e({open_n23283,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c6_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c6_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c6_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c6_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c6_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c6_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c6_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c6_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c6_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c6_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c6_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c6_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_025 ,\picorv32_core/cpuregs_p2/dram_do_i1_024 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c6_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c6_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c6_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c6_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c6_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c6_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c6_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_027 ,\picorv32_core/cpuregs_p2/dram_do_i1_026 }));
  EG_PHY_LSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c7_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \picorv32_core/cpuregs_p2/dram_r1_c7_l  (
    .a({\picorv32_core/cpuregs_wrdata [28],\picorv32_core/latched_rd [0]}),
    .b({\picorv32_core/cpuregs_wrdata [29],\picorv32_core/latched_rd [1]}),
    .c({\picorv32_core/cpuregs_wrdata [30],\picorv32_core/latched_rd [2]}),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_wrdata [31],\picorv32_core/latched_rd [3]}),
    .e({open_n23318,\picorv32_core/n456_1_al_n604 }),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c7_di ),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c7_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c7_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c7_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c7_we ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c7_l"),
    //.R_POSITION("X0Y0Z0"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c7_m0  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c7_di [1:0]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c7_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c7_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c7_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c7_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_029 ,\picorv32_core/cpuregs_p2/dram_do_i1_028 }));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/cpuregs_p2/dram_r1_c7_l"),
    //.R_POSITION("X0Y0Z1"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"))
    \picorv32_core/cpuregs_p2/dram_r1_c7_m1  (
    .a({\picorv32_core/decoded_rs2 [0],\picorv32_core/decoded_rs2 [0]}),
    .b({\picorv32_core/decoded_rs2 [1],\picorv32_core/decoded_rs2 [1]}),
    .c({\picorv32_core/decoded_rs2 [2],\picorv32_core/decoded_rs2 [2]}),
    .d({\picorv32_core/decoded_rs2 [3],\picorv32_core/decoded_rs2 [3]}),
    .dpram_di(\picorv32_core/cpuregs_p2/dram_r1_c7_di [3:2]),
    .dpram_mode(\picorv32_core/cpuregs_p2/dram_r1_c7_mode ),
    .dpram_waddr(\picorv32_core/cpuregs_p2/dram_r1_c7_waddr ),
    .dpram_wclk(\picorv32_core/cpuregs_p2/dram_r1_c7_wclk ),
    .dpram_we(\picorv32_core/cpuregs_p2/dram_r1_c7_we ),
    .f({\picorv32_core/cpuregs_p2/dram_do_i1_031 ,\picorv32_core/cpuregs_p2/dram_do_i1_030 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*C*~(A*~(B*D)))"),
    //.LUT1("(~1*C*~(A*~(B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101000001010000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/decoder_pseudo_trigger_reg  (
    .a({_al_u1088_o,_al_u1088_o}),
    .b({\picorv32_core/mem_xfer_placeOpt_1 ,\picorv32_core/mem_xfer_placeOpt_1 }),
    .c({\picorv32_core/n16 ,\picorv32_core/n16 }),
    .clk(clk_pad),
    .d({\picorv32_core/n180 ,\picorv32_core/n180 }),
    .mi({open_n23363,\picorv32_core/mem_do_prefetch }),
    .sr(\picorv32_core/u625_sel_is_2_o ),
    .fx({open_n23367,\picorv32_core/n580 }),
    .q({open_n23368,\picorv32_core/decoder_pseudo_trigger }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~(~A*~B)*~(0*~C)))"),
    //.LUT1("(D*~(~(~B*~A)*~(1*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100000000),
    .INIT_LUT1(16'b0001111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/decoder_trigger_reg  (
    .a({_al_u1184_o,\picorv32_core/mem_do_prefetch }),
    .b({\picorv32_core/mem_do_prefetch ,_al_u1184_o}),
    .c({_al_u1906_o,_al_u1906_o}),
    .clk(clk_pad),
    .d({_al_u1546_o,_al_u1546_o}),
    .mi({open_n23380,\picorv32_core/mem_do_rinst }),
    .q({open_n23387,\picorv32_core/decoder_trigger }));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(~D*~C*~A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/instr_add_reg|picorv32_core/instr_sltu_reg  (
    .a({\picorv32_core/mem_rdata_q [12],_al_u976_o}),
    .b({_al_u976_o,\picorv32_core/mem_rdata_q [12]}),
    .c({\picorv32_core/mem_rdata_q [13],\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [14],\picorv32_core/mem_rdata_q [14]}),
    .sr(resetn_placeOpt_8),
    .q({\picorv32_core/instr_add ,\picorv32_core/instr_sltu }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/instr_addi_reg|picorv32_core/instr_sltiu_reg  (
    .a({\picorv32_core/is_alu_reg_imm ,\picorv32_core/is_alu_reg_imm }),
    .b({\picorv32_core/mem_rdata_q [12],\picorv32_core/mem_rdata_q [12]}),
    .c({\picorv32_core/mem_rdata_q [13],\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [14],\picorv32_core/mem_rdata_q [14]}),
    .sr(resetn_placeOpt_8),
    .q({\picorv32_core/instr_addi ,\picorv32_core/instr_sltiu }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/instr_and_reg|picorv32_core/instr_xor_reg  (
    .a({_al_u976_o,_al_u976_o}),
    .b({\picorv32_core/mem_rdata_q [12],\picorv32_core/mem_rdata_q [12]}),
    .c({\picorv32_core/mem_rdata_q [13],\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [14],\picorv32_core/mem_rdata_q [14]}),
    .sr(resetn_placeOpt_8),
    .q({\picorv32_core/instr_and ,\picorv32_core/instr_xor }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/instr_beq_reg|picorv32_core/instr_bltu_reg  (
    .a({\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ,\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .b({\picorv32_core/mem_rdata_q [12],\picorv32_core/mem_rdata_q [12]}),
    .c({\picorv32_core/mem_rdata_q [13],\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [14],\picorv32_core/mem_rdata_q [14]}),
    .sr(resetn_placeOpt_8),
    .q({\picorv32_core/instr_beq ,\picorv32_core/instr_bltu }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(0*C*A))"),
    //.LUT1("~(~(D*B)*~(1*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110000000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/instr_jal_reg  (
    .a({_al_u1535_o,_al_u1535_o}),
    .b({_al_u1536_o,_al_u1536_o}),
    .c({_al_u1533_o,_al_u1533_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mux81_sel_is_1_o ,\picorv32_core/mux81_sel_is_1_o }),
    .mi({open_n23466,\picorv32_core/mem_rdata_latched [3]}),
    .q({open_n23473,\picorv32_core/instr_jal }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("A*B*~C*~D+A*B*C*~D"),
    //.LUTF1("0"),
    //.LUTG0("0"),
    //.LUTG1("~D*~B*~A*~C+~D*~B*~A*C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010001000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/instr_lb_reg|picorv32_core/instr_lh_reg  (
    .a({\picorv32_core/mem_rdata_q [13],\picorv32_core/is_lb_lh_lw_lbu_lhu }),
    .b({\picorv32_core/mem_rdata_q [12],\picorv32_core/mem_rdata_q [12]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [14],\picorv32_core/mem_rdata_q [14]}),
    .e({\picorv32_core/is_lb_lh_lw_lbu_lhu ,\picorv32_core/mem_rdata_q [13]}),
    .q({\picorv32_core/instr_lb ,\picorv32_core/instr_lh }));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~C*~B*~(A*~D))"),
    //.LUTF1("0"),
    //.LUTG0("(~1*~C*~B*~(A*~D))"),
    //.LUTG1("D*~A*~C*~B+D*~A*~C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000001),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/instr_lbu_reg|_al_u1908  (
    .a({\picorv32_core/mem_rdata_q [12],\picorv32_core/mem_do_prefetch_placeOpt_8 }),
    .b({open_n23496,\picorv32_core/instr_lb }),
    .c({\picorv32_core/mem_rdata_q [13],\picorv32_core/instr_lbu }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [14],_al_u1546_o}),
    .e({\picorv32_core/is_lb_lh_lw_lbu_lhu ,\picorv32_core/mem_do_rdata }),
    .f({open_n23512,_al_u1908_o}),
    .q({\picorv32_core/instr_lbu ,open_n23516}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*A)"),
    //.LUTF1("0"),
    //.LUTG0("(D*~C*B*A)"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/instr_lw_reg|picorv32_core/instr_lhu_reg  (
    .a({\picorv32_core/n289_lutinv ,\picorv32_core/is_lb_lh_lw_lbu_lhu }),
    .b({open_n23517,\picorv32_core/mem_rdata_q [12]}),
    .c({open_n23518,\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({open_n23519,\picorv32_core/mem_rdata_q [14]}),
    .e({\picorv32_core/is_lb_lh_lw_lbu_lhu ,open_n23520}),
    .q({\picorv32_core/instr_lw ,\picorv32_core/instr_lhu }));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*B*A)"),
    //.LUTF1("0"),
    //.LUTG0("(1*D*~C*B*A)"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/instr_rdcycleh_reg|_al_u1098  (
    .a({_al_u1098_o,_al_u1097_o}),
    .b({open_n23541,\picorv32_core/mem_rdata_q [27]}),
    .c({open_n23542,\picorv32_core/mem_rdata_q [29]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({open_n23543,\picorv32_core/mem_rdata_q [30]}),
    .e({_al_u1143_o,\picorv32_core/mem_rdata_q [31]}),
    .f({open_n23559,_al_u1098_o}),
    .q({\picorv32_core/instr_rdcycleh ,open_n23563}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/instr_rdinstr_reg|picorv32_core/instr_rdinstrh_reg  (
    .b({_al_u1100_o,open_n23566}),
    .c({open_n23567,_al_u1098_o}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .e({_al_u1095_o,_al_u1095_o}),
    .q({\picorv32_core/instr_rdinstr ,\picorv32_core/instr_rdinstrh }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*C*B*A)"),
    //.LUT1("(~1*~D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/instr_slli_reg  (
    .a({\picorv32_core/n304_lutinv ,\picorv32_core/n304_lutinv }),
    .b({\picorv32_core/is_alu_reg_imm ,\picorv32_core/is_alu_reg_imm }),
    .c({\picorv32_core/mem_rdata_q [12],\picorv32_core/mem_rdata_q [12]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [13],\picorv32_core/mem_rdata_q [13]}),
    .mi({open_n23600,\picorv32_core/mem_rdata_q [14]}),
    .q({open_n23607,\picorv32_core/instr_slli }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("0"),
    //.LUTG0("A*~D*B*~C+A*~D*B*C"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000010001000),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/instr_slt_reg|picorv32_core/instr_or_reg  (
    .a({open_n23608,_al_u976_o}),
    .b({_al_u976_o,\picorv32_core/mem_rdata_q [13]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({open_n23611,\picorv32_core/mem_rdata_q [12]}),
    .e({\picorv32_core/n289_lutinv ,\picorv32_core/mem_rdata_q [14]}),
    .sr(resetn_placeOpt_8),
    .q({\picorv32_core/instr_slt ,\picorv32_core/instr_or }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~D*C*B*A)"),
    //.LUT1("(1*~D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000010000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/instr_srli_reg  (
    .a({\picorv32_core/n304_lutinv ,\picorv32_core/n304_lutinv }),
    .b({\picorv32_core/is_alu_reg_imm ,\picorv32_core/is_alu_reg_imm }),
    .c({\picorv32_core/mem_rdata_q [12],\picorv32_core/mem_rdata_q [12]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [13],\picorv32_core/mem_rdata_q [13]}),
    .mi({open_n23641,\picorv32_core/mem_rdata_q [14]}),
    .q({open_n23648,\picorv32_core/instr_srli }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(~B*A*~(0*D)))"),
    //.LUT1("~(~C*~(~B*A*~(1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001011110010),
    .INIT_LUT1(16'b1111000011110010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/is_alu_reg_imm_reg  (
    .a({_al_u1649_o,_al_u1649_o}),
    .b({_al_u1653_o,_al_u1653_o}),
    .c({_al_u1652_o,_al_u1652_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u1651_o,_al_u1651_o}),
    .mi({open_n23659,_al_u1654_o}),
    .q({open_n23666,\picorv32_core/is_alu_reg_imm }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D*~(0*A*~B))"),
    //.LUT1("~(~C*~D*~(1*A*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111111111110010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/is_alu_reg_reg_reg  (
    .a({\picorv32_core/n98_lutinv ,\picorv32_core/n98_lutinv }),
    .b({_al_u1605_o,_al_u1605_o}),
    .c({_al_u1604_o,_al_u1604_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u1603_o,_al_u1603_o}),
    .mi({open_n23677,_al_u1606_o}),
    .q({open_n23684,\picorv32_core/is_alu_reg_reg }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~D*~C*~B*~A)"),
    //.LUT1("~(~1*~B*~C*~D*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111110),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/is_compare_reg  (
    .a({\picorv32_core/instr_slt ,\picorv32_core/instr_slt }),
    .b({\picorv32_core/instr_sltu ,\picorv32_core/instr_slti }),
    .c({\picorv32_core/instr_sltiu ,\picorv32_core/instr_sltiu }),
    .clk(clk_pad),
    .d({\picorv32_core/instr_slti ,\picorv32_core/instr_sltu }),
    .mi({open_n23696,\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .sr(\picorv32_core/u449_sel_is_0_o ),
    .q({open_n23702,\picorv32_core/is_compare }));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(~0*~A*B)*~(C*D))"),
    //.LUT1("~(~(~1*~B*C)*~(A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010001000100),
    .INIT_LUT1(16'b1010101000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/is_lb_lh_lw_lbu_lhu_reg  (
    .a({_al_u1593_o,\picorv32_core/mem_rdata_latched$0$_placeOpt_1 }),
    .b({\picorv32_core/mem_rdata_latched$0$_placeOpt_1 ,_al_u1597_o}),
    .c({_al_u1597_o,_al_u1593_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u1596_o,_al_u1596_o}),
    .mi({open_n23713,_al_u1481_o_placeOpt_3}),
    .q({open_n23720,\picorv32_core/is_lb_lh_lw_lbu_lhu }));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~C*~B*~(A*~D))"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~1*~C*~B*~(A*~D))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000001),
    .INIT_LUTF1(16'b1111111110101010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/is_lbu_lhu_lw_reg|_al_u1914  (
    .a({\picorv32_core/instr_lw ,\picorv32_core/mem_do_prefetch_placeOpt_5 }),
    .b({open_n23721,\picorv32_core/instr_lh }),
    .c({open_n23722,\picorv32_core/instr_lhu }),
    .clk(clk_pad),
    .d({\picorv32_core/instr_lhu ,_al_u1546_o_placeOpt_8}),
    .e({\picorv32_core/instr_lbu ,\picorv32_core/mem_do_rdata }),
    .f({\picorv32_core/n168 ,_al_u1914_o}),
    .q({\picorv32_core/is_lbu_lhu_lw ,open_n23742}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~C*~A*~B*~D)"),
    //.LUT1("~(~1*~C*~A*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111110),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub_reg  (
    .a({\picorv32_core/instr_addi ,\picorv32_core/instr_addi }),
    .b({\picorv32_core/instr_add ,\picorv32_core/instr_add }),
    .c({\picorv32_core/instr_jalr ,\picorv32_core/instr_jalr }),
    .clk(clk_pad),
    .d({\picorv32_core/n472 ,\picorv32_core/n472 }),
    .mi({open_n23754,\picorv32_core/instr_sub }),
    .sr(\picorv32_core/n274 ),
    .fx({open_n23758,\picorv32_core/n165 }),
    .q({open_n23759,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/is_sll_srl_sra_reg|picorv32_core/is_slli_srli_srai_reg  (
    .c({\picorv32_core/is_alu_reg_reg ,\picorv32_core/is_alu_reg_imm }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({_al_u1102_o,_al_u1102_o}),
    .q({\picorv32_core/is_sll_srl_sra ,\picorv32_core/is_slli_srli_srai }));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("C*~D*~A*~B+C*~D*A*~B+C*~D*~A*B"),
    //.LUTF1("~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*B*~D*C+A*B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG0("C*~D*A*~B"),
    //.LUTG1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000001110000),
    .INIT_LUTF1(16'b1111111111001100),
    .INIT_LUTG0(16'b0000000000100000),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/is_slti_blt_slt_reg|_al_u1215  (
    .a({open_n23782,\picorv32_core/alu_lts }),
    .b({\picorv32_core/instr_slti ,\picorv32_core/is_slti_blt_slt }),
    .c({open_n23783,_al_u1213_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_slt ,_al_u1214_o}),
    .e({\picorv32_core/instr_blt ,\picorv32_core/instr_bge }),
    .f({open_n23800,_al_u1215_o}),
    .q({\picorv32_core/is_slti_blt_slt ,open_n23804}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~D*~C+A*~B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~B*~D*~C+A*~B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*~B*D*C+A*~B*D*C"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100110011),
    .INIT_LUTF1(16'b1111110011111100),
    .INIT_LUTG0(16'b0011001100110011),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/is_sltiu_bltu_sltu_reg|picorv32_core/reg14_b0  (
    .b({\picorv32_core/instr_sltiu ,_al_u1293_o}),
    .c({\picorv32_core/instr_sltu ,open_n23807}),
    .clk(clk_pad),
    .d({open_n23809,\picorv32_core/is_compare }),
    .e({\picorv32_core/instr_bltu ,_al_u1216_o}),
    .q({\picorv32_core/is_sltiu_bltu_sltu ,\picorv32_core/alu_out_q [0]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~(~A*~(D)*~(0)+~A*D*~(0)+~(~A)*D*0+~A*D*0)))"),
    //.LUT1("~(B*~(A*~(~C*~(D)*~(1)+~C*D*~(1)+~(~C)*D*1+~C*D*1)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011001110110011),
    .INIT_LUT1(16'b0011001110111011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/latched_branch_reg  (
    .a({\picorv32_core/n666_lutinv ,\picorv32_core/instr_jalr }),
    .b({_al_u1285_o,_al_u1285_o}),
    .c({\picorv32_core/instr_jalr ,\picorv32_core/n666_lutinv }),
    .clk(clk_pad),
    .d({_al_u1216_o,_al_u1216_o}),
    .mi({open_n23841,\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .sr(resetn_placeOpt_10),
    .q({open_n23847,\picorv32_core/latched_branch }));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*C*A*~(0)+D*B*C*A*~(0)+~(D)*~(B)*~(C)*~(A)*0+D*~(B)*~(C)*~(A)*0+~(D)*~(B)*C*~(A)*0+D*~(B)*C*~(A)*0+~(D)*B*C*~(A)*0+~(D)*~(B)*~(C)*A*0+D*~(B)*~(C)*A*0+~(D)*~(B)*C*A*0+D*~(B)*C*A*0+~(D)*B*C*A*0+D*B*C*A*0)"),
    //.LUTF1("(D*~(C)*B*A*~(0)+D*C*B*A*~(0)+~(D)*~(C)*~(B)*~(A)*0+D*~(C)*~(B)*~(A)*0+~(D)*~(C)*B*~(A)*0+D*~(C)*B*~(A)*0+~(D)*C*B*~(A)*0+~(D)*~(C)*~(B)*A*0+D*~(C)*~(B)*A*0+~(D)*~(C)*B*A*0+D*~(C)*B*A*0+~(D)*C*B*A*0+D*C*B*A*0)"),
    //.LUTG0("(D*~(B)*C*A*~(1)+D*B*C*A*~(1)+~(D)*~(B)*~(C)*~(A)*1+D*~(B)*~(C)*~(A)*1+~(D)*~(B)*C*~(A)*1+D*~(B)*C*~(A)*1+~(D)*B*C*~(A)*1+~(D)*~(B)*~(C)*A*1+D*~(B)*~(C)*A*1+~(D)*~(B)*C*A*1+D*~(B)*C*A*1+~(D)*B*C*A*1+D*B*C*A*1)"),
    //.LUTG1("(D*~(C)*B*A*~(1)+D*C*B*A*~(1)+~(D)*~(C)*~(B)*~(A)*1+D*~(C)*~(B)*~(A)*1+~(D)*~(C)*B*~(A)*1+D*~(C)*B*~(A)*1+~(D)*C*B*~(A)*1+~(D)*~(C)*~(B)*A*1+D*~(C)*~(B)*A*1+~(D)*~(C)*B*A*1+D*~(C)*B*A*1+~(D)*C*B*A*1+D*C*B*A*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010000000000000),
    .INIT_LUTF1(16'b1000100000000000),
    .INIT_LUTG0(16'b1011001111110011),
    .INIT_LUTG1(16'b1000111111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/latched_is_lh_reg|picorv32_core/latched_is_lb_reg  (
    .a({\picorv32_core/instr_lh ,\picorv32_core/instr_lb }),
    .b({\picorv32_core/n669_lutinv_placeOpt_4 ,_al_u1609_o}),
    .c({_al_u1609_o,\picorv32_core/n669_lutinv_placeOpt_4 }),
    .clk(clk_pad),
    .d({\picorv32_core/mux132_b0_sel_is_3_o ,\picorv32_core/mux132_b0_sel_is_3_o }),
    .e({\picorv32_core/latched_is_lh ,\picorv32_core/latched_is_lb }),
    .sr(resetn_placeOpt_17),
    .q({\picorv32_core/latched_is_lh ,\picorv32_core/latched_is_lb }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*C*A*~(0)+D*B*C*A*~(0)+~(D)*~(B)*~(C)*~(A)*0+D*~(B)*~(C)*~(A)*0+~(D)*~(B)*C*~(A)*0+D*~(B)*C*~(A)*0+~(D)*B*C*~(A)*0+~(D)*~(B)*~(C)*A*0+D*~(B)*~(C)*A*0+~(D)*~(B)*C*A*0+D*~(B)*C*A*0+~(D)*B*C*A*0+D*B*C*A*0)"),
    //.LUT1("(D*~(B)*C*A*~(1)+D*B*C*A*~(1)+~(D)*~(B)*~(C)*~(A)*1+D*~(B)*~(C)*~(A)*1+~(D)*~(B)*C*~(A)*1+D*~(B)*C*~(A)*1+~(D)*B*C*~(A)*1+~(D)*~(B)*~(C)*A*1+D*~(B)*~(C)*A*1+~(D)*~(B)*C*A*1+D*~(B)*C*A*1+~(D)*B*C*A*1+D*B*C*A*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010000000000000),
    .INIT_LUT1(16'b1011001111110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/latched_is_lu_reg  (
    .a({\picorv32_core/is_lbu_lhu_lw ,\picorv32_core/is_lbu_lhu_lw }),
    .b({_al_u1609_o,_al_u1609_o}),
    .c({\picorv32_core/n669_lutinv_placeOpt_4 ,\picorv32_core/n669_lutinv_placeOpt_4 }),
    .clk(clk_pad),
    .d({\picorv32_core/mux132_b0_sel_is_3_o ,\picorv32_core/mux132_b0_sel_is_3_o }),
    .mi({open_n23879,\picorv32_core/latched_is_lu }),
    .sr(resetn_placeOpt_17),
    .q({open_n23885,\picorv32_core/latched_is_lu }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_0|picorv32_core/lt0_cin  (
    .a({\picorv32_core/pcpi_rs1$0$ ,1'b0}),
    .b({mem_la_wdata[0],open_n23886}),
    .fco(\picorv32_core/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_10|picorv32_core/lt0_9  (
    .a({\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$9$ }),
    .b({\picorv32_core/pcpi_rs2$10$ ,\picorv32_core/pcpi_rs2$9$ }),
    .fci(\picorv32_core/lt0_c9 ),
    .fco(\picorv32_core/lt0_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_12|picorv32_core/lt0_11  (
    .a({\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/pcpi_rs1$11$ }),
    .b({\picorv32_core/pcpi_rs2$12$ ,\picorv32_core/pcpi_rs2$11$ }),
    .fci(\picorv32_core/lt0_c11 ),
    .fco(\picorv32_core/lt0_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_14|picorv32_core/lt0_13  (
    .a({\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$13$ }),
    .b({\picorv32_core/pcpi_rs2$14$ ,\picorv32_core/pcpi_rs2$13$ }),
    .fci(\picorv32_core/lt0_c13 ),
    .fco(\picorv32_core/lt0_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_16|picorv32_core/lt0_15  (
    .a({\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/pcpi_rs1$15$ }),
    .b({\picorv32_core/pcpi_rs2$16$ ,\picorv32_core/pcpi_rs2$15$ }),
    .fci(\picorv32_core/lt0_c15 ),
    .fco(\picorv32_core/lt0_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_18|picorv32_core/lt0_17  (
    .a({\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$17$ }),
    .b({\picorv32_core/pcpi_rs2$18$ ,\picorv32_core/pcpi_rs2$17$ }),
    .fci(\picorv32_core/lt0_c17 ),
    .fco(\picorv32_core/lt0_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_20|picorv32_core/lt0_19  (
    .a({\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/pcpi_rs1$19$ }),
    .b({\picorv32_core/pcpi_rs2$20$ ,\picorv32_core/pcpi_rs2$19$ }),
    .fci(\picorv32_core/lt0_c19 ),
    .fco(\picorv32_core/lt0_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_22|picorv32_core/lt0_21  (
    .a({\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs1$21$ }),
    .b({\picorv32_core/pcpi_rs2$22$ ,\picorv32_core/pcpi_rs2$21$ }),
    .fci(\picorv32_core/lt0_c21 ),
    .fco(\picorv32_core/lt0_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_24|picorv32_core/lt0_23  (
    .a({\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/pcpi_rs1$23$ }),
    .b({\picorv32_core/pcpi_rs2$24$ ,\picorv32_core/pcpi_rs2$23$ }),
    .fci(\picorv32_core/lt0_c23 ),
    .fco(\picorv32_core/lt0_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_26|picorv32_core/lt0_25  (
    .a({\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$25$ }),
    .b({\picorv32_core/pcpi_rs2$26$ ,\picorv32_core/pcpi_rs2$25$ }),
    .fci(\picorv32_core/lt0_c25 ),
    .fco(\picorv32_core/lt0_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_28|picorv32_core/lt0_27  (
    .a({\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/pcpi_rs1$27$ }),
    .b({\picorv32_core/pcpi_rs2$28$ ,\picorv32_core/pcpi_rs2$27$ }),
    .fci(\picorv32_core/lt0_c27 ),
    .fco(\picorv32_core/lt0_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_2|picorv32_core/lt0_1  (
    .a({\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$1$ }),
    .b(mem_la_wdata[2:1]),
    .fci(\picorv32_core/lt0_c1 ),
    .fco(\picorv32_core/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_30|picorv32_core/lt0_29  (
    .a({\picorv32_core/pcpi_rs1$30$ ,\picorv32_core/pcpi_rs1$29$ }),
    .b({\picorv32_core/pcpi_rs2$30$ ,\picorv32_core/pcpi_rs2$29$ }),
    .fci(\picorv32_core/lt0_c29 ),
    .fco(\picorv32_core/lt0_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_4|picorv32_core/lt0_3  (
    .a({\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/pcpi_rs1$3$ }),
    .b(mem_la_wdata[4:3]),
    .fci(\picorv32_core/lt0_c3 ),
    .fco(\picorv32_core/lt0_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_6|picorv32_core/lt0_5  (
    .a({\picorv32_core/pcpi_rs1$6$ ,\picorv32_core/pcpi_rs1$5$ }),
    .b(mem_la_wdata[6:5]),
    .fci(\picorv32_core/lt0_c5 ),
    .fco(\picorv32_core/lt0_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_8|picorv32_core/lt0_7  (
    .a({\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/pcpi_rs1$7$ }),
    .b({\picorv32_core/pcpi_rs2$8$ ,mem_la_wdata[7]}),
    .fci(\picorv32_core/lt0_c7 ),
    .fco(\picorv32_core/lt0_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt0_0|picorv32_core/lt0_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt0_cout|picorv32_core/lt0_31  (
    .a({1'b0,\picorv32_core/pcpi_rs2$31$ }),
    .b({1'b1,\picorv32_core/pcpi_rs1$31$ }),
    .fci(\picorv32_core/lt0_c31 ),
    .f({\picorv32_core/alu_lts ,open_n24290}));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_0|picorv32_core/lt1_cin  (
    .a({\picorv32_core/pcpi_rs1$0$ ,1'b0}),
    .b({mem_la_wdata[0],open_n24296}),
    .fco(\picorv32_core/lt1_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_10|picorv32_core/lt1_9  (
    .a({\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$9$ }),
    .b({\picorv32_core/pcpi_rs2$10$ ,\picorv32_core/pcpi_rs2$9$ }),
    .fci(\picorv32_core/lt1_c9 ),
    .fco(\picorv32_core/lt1_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_12|picorv32_core/lt1_11  (
    .a({\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/pcpi_rs1$11$ }),
    .b({\picorv32_core/pcpi_rs2$12$ ,\picorv32_core/pcpi_rs2$11$ }),
    .fci(\picorv32_core/lt1_c11 ),
    .fco(\picorv32_core/lt1_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_14|picorv32_core/lt1_13  (
    .a({\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$13$ }),
    .b({\picorv32_core/pcpi_rs2$14$ ,\picorv32_core/pcpi_rs2$13$ }),
    .fci(\picorv32_core/lt1_c13 ),
    .fco(\picorv32_core/lt1_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_16|picorv32_core/lt1_15  (
    .a({\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/pcpi_rs1$15$ }),
    .b({\picorv32_core/pcpi_rs2$16$ ,\picorv32_core/pcpi_rs2$15$ }),
    .fci(\picorv32_core/lt1_c15 ),
    .fco(\picorv32_core/lt1_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_18|picorv32_core/lt1_17  (
    .a({\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$17$ }),
    .b({\picorv32_core/pcpi_rs2$18$ ,\picorv32_core/pcpi_rs2$17$ }),
    .fci(\picorv32_core/lt1_c17 ),
    .fco(\picorv32_core/lt1_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_20|picorv32_core/lt1_19  (
    .a({\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/pcpi_rs1$19$ }),
    .b({\picorv32_core/pcpi_rs2$20$ ,\picorv32_core/pcpi_rs2$19$ }),
    .fci(\picorv32_core/lt1_c19 ),
    .fco(\picorv32_core/lt1_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_22|picorv32_core/lt1_21  (
    .a({\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs1$21$ }),
    .b({\picorv32_core/pcpi_rs2$22$ ,\picorv32_core/pcpi_rs2$21$ }),
    .fci(\picorv32_core/lt1_c21 ),
    .fco(\picorv32_core/lt1_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_24|picorv32_core/lt1_23  (
    .a({\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/pcpi_rs1$23$ }),
    .b({\picorv32_core/pcpi_rs2$24$ ,\picorv32_core/pcpi_rs2$23$ }),
    .fci(\picorv32_core/lt1_c23 ),
    .fco(\picorv32_core/lt1_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_26|picorv32_core/lt1_25  (
    .a({\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$25$ }),
    .b({\picorv32_core/pcpi_rs2$26$ ,\picorv32_core/pcpi_rs2$25$ }),
    .fci(\picorv32_core/lt1_c25 ),
    .fco(\picorv32_core/lt1_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_28|picorv32_core/lt1_27  (
    .a({\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/pcpi_rs1$27$ }),
    .b({\picorv32_core/pcpi_rs2$28$ ,\picorv32_core/pcpi_rs2$27$ }),
    .fci(\picorv32_core/lt1_c27 ),
    .fco(\picorv32_core/lt1_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_2|picorv32_core/lt1_1  (
    .a({\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$1$ }),
    .b(mem_la_wdata[2:1]),
    .fci(\picorv32_core/lt1_c1 ),
    .fco(\picorv32_core/lt1_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_30|picorv32_core/lt1_29  (
    .a({\picorv32_core/pcpi_rs1$30$ ,\picorv32_core/pcpi_rs1$29$ }),
    .b({\picorv32_core/pcpi_rs2$30$ ,\picorv32_core/pcpi_rs2$29$ }),
    .fci(\picorv32_core/lt1_c29 ),
    .fco(\picorv32_core/lt1_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_4|picorv32_core/lt1_3  (
    .a({\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/pcpi_rs1$3$ }),
    .b(mem_la_wdata[4:3]),
    .fci(\picorv32_core/lt1_c3 ),
    .fco(\picorv32_core/lt1_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_6|picorv32_core/lt1_5  (
    .a({\picorv32_core/pcpi_rs1$6$ ,\picorv32_core/pcpi_rs1$5$ }),
    .b(mem_la_wdata[6:5]),
    .fci(\picorv32_core/lt1_c5 ),
    .fco(\picorv32_core/lt1_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_8|picorv32_core/lt1_7  (
    .a({\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/pcpi_rs1$7$ }),
    .b({\picorv32_core/pcpi_rs2$8$ ,mem_la_wdata[7]}),
    .fci(\picorv32_core/lt1_c7 ),
    .fco(\picorv32_core/lt1_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt1_0|picorv32_core/lt1_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt1_cout|picorv32_core/lt1_31  (
    .a({1'b0,\picorv32_core/pcpi_rs1$31$ }),
    .b({1'b1,\picorv32_core/pcpi_rs2$31$ }),
    .fci(\picorv32_core/lt1_c31 ),
    .f({\picorv32_core/alu_ltu ,open_n24700}));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt2_0|picorv32_core/lt2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt2_0|picorv32_core/lt2_cin  (
    .a(2'b01),
    .b({\picorv32_core/reg_sh [0],open_n24706}),
    .fco(\picorv32_core/lt2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt2_0|picorv32_core/lt2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt2_2|picorv32_core/lt2_1  (
    .a(2'b10),
    .b(\picorv32_core/reg_sh [2:1]),
    .fci(\picorv32_core/lt2_c1 ),
    .fco(\picorv32_core/lt2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt2_0|picorv32_core/lt2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt2_4|picorv32_core/lt2_3  (
    .a(2'b00),
    .b(\picorv32_core/reg_sh [4:3]),
    .fci(\picorv32_core/lt2_c3 ),
    .fco(\picorv32_core/lt2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/lt2_0|picorv32_core/lt2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \picorv32_core/lt2_cout_al_u2576  (
    .a({open_n24780,1'b0}),
    .b({open_n24781,1'b1}),
    .fci(\picorv32_core/lt2_c5 ),
    .f({open_n24800,\picorv32_core/n554 }));
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))*~(A)+~0*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*~(A)+~(~0)*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A+~0*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A)"),
    //.LUT1("~(~1*~((~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))*~(A)+~1*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*~(A)+~(~1)*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A+~1*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010101000001000),
    .INIT_LUT1(16'b0111111101011101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b0  (
    .a({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({_al_u1088_o,_al_u1088_o}),
    .c({_al_u1282_o,_al_u1282_o}),
    .ce(\picorv32_core/mem_xfer_placeOpt_3 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched_noshuffle [0],\picorv32_core/mem_rdata_latched_noshuffle [0]}),
    .mi({open_n24816,\picorv32_core/mem_16bit_buffer [0]}),
    .fx({open_n24821,\picorv32_core/mem_rdata_latched [0]}),
    .q({open_n24822,\picorv32_core/mem_rdata_q [0]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))*~(C)+~0*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*~(C)+~(~0)*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C+~0*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C)"),
    //.LUT1("~(~1*~((~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))*~(C)+~1*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*~(C)+~(~1)*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C+~1*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000011100000),
    .INIT_LUT1(16'b0010111111101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b0_placeOpt_1  (
    .a({\picorv32_core/mem_rdata_latched_noshuffle [0],\picorv32_core/mem_rdata_latched_noshuffle [0]}),
    .b({_al_u1088_o,_al_u1088_o}),
    .c({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .ce(\picorv32_core/mem_xfer_placeOpt_3 ),
    .clk(clk_pad),
    .d({_al_u1282_o,_al_u1282_o}),
    .mi({open_n24833,\picorv32_core/mem_16bit_buffer [0]}),
    .fx({open_n24838,\picorv32_core/mem_rdata_latched$0$_placeOpt_1 }));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))*~(C)+~0*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*~(C)+~(~0)*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C+~0*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C)"),
    //.LUT1("~(~1*~((~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))*~(C)+~1*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*~(C)+~(~1)*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C+~1*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000011100000),
    .INIT_LUT1(16'b0010111111101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b0_placeOpt_2  (
    .a({\picorv32_core/mem_rdata_latched_noshuffle [0],\picorv32_core/mem_rdata_latched_noshuffle [0]}),
    .b({_al_u1088_o,_al_u1088_o}),
    .c({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .ce(\picorv32_core/mem_xfer_placeOpt_3 ),
    .clk(clk_pad),
    .d({_al_u1282_o,_al_u1282_o}),
    .mi({open_n24851,\picorv32_core/mem_16bit_buffer [0]}),
    .fx({open_n24856,\picorv32_core/mem_rdata_latched$0$_placeOpt_2 }));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))*~(A)+~0*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*~(A)+~(~0)*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A+~0*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A)"),
    //.LUT1("~(~1*~((~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))*~(B)+~1*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*~(B)+~(~1)*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B+~1*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010101000001000),
    .INIT_LUT1(16'b0111111100111011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b0_placeOpt_3  (
    .a({_al_u1088_o,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,_al_u1088_o}),
    .c({_al_u1282_o,_al_u1282_o}),
    .ce(\picorv32_core/mem_xfer_placeOpt_3 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched_noshuffle [0],\picorv32_core/mem_rdata_latched_noshuffle [0]}),
    .mi({open_n24869,\picorv32_core/mem_16bit_buffer [0]}),
    .fx({open_n24874,\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))*~(C)+~0*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*~(C)+~(~0)*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C+~0*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C)"),
    //.LUT1("~(~1*~((~B*~(D)*~(A)+~B*D*~(A)+~(~B)*D*A+~B*D*A))*~(C)+~1*(~B*~(D)*~(A)+~B*D*~(A)+~(~B)*D*A+~B*D*A)*~(C)+~(~1)*(~B*~(D)*~(A)+~B*D*~(A)+~(~B)*D*A+~B*D*A)*C+~1*(~B*~(D)*~(A)+~B*D*~(A)+~(~B)*D*A+~B*D*A)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000011100000),
    .INIT_LUT1(16'b0100111111101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b0_placeOpt_4  (
    .a({_al_u1088_o,\picorv32_core/mem_rdata_latched_noshuffle [0]}),
    .b({\picorv32_core/mem_rdata_latched_noshuffle [0],_al_u1088_o}),
    .c({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .ce(\picorv32_core/mem_xfer_placeOpt_3 ),
    .clk(clk_pad),
    .d({_al_u1282_o,_al_u1282_o}),
    .mi({open_n24887,\picorv32_core/mem_16bit_buffer [0]}),
    .fx({open_n24892,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))*~(C)+~0*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*~(C)+~(~0)*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C+~0*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C)"),
    //.LUT1("~(~1*~((~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))*~(C)+~1*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*~(C)+~(~1)*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C+~1*(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000011100000),
    .INIT_LUT1(16'b0010111111101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b0_placeOpt_5  (
    .a({\picorv32_core/mem_rdata_latched_noshuffle [0],\picorv32_core/mem_rdata_latched_noshuffle [0]}),
    .b({_al_u1088_o,_al_u1088_o}),
    .c({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .ce(\picorv32_core/mem_xfer_placeOpt_3 ),
    .clk(clk_pad),
    .d({_al_u1282_o,_al_u1282_o}),
    .mi({open_n24905,\picorv32_core/mem_16bit_buffer [0]}),
    .fx({open_n24910,\picorv32_core/mem_rdata_latched$0$_placeOpt_5 }));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))*~(B)+~0*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*~(B)+~(~0)*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B+~0*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B)"),
    //.LUT1("~(~1*~((~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))*~(A)+~1*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*~(A)+~(~1)*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A+~1*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100110000001000),
    .INIT_LUT1(16'b0111111101011101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b1  (
    .a({\picorv32_core/mux4_b0_sel_is_0_o ,_al_u1088_o}),
    .b({_al_u1088_o,\picorv32_core/mux4_b0_sel_is_0_o }),
    .c({_al_u1276_o,_al_u1276_o}),
    .ce(\picorv32_core/mem_xfer_placeOpt_3 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched_noshuffle [1],\picorv32_core/mem_rdata_latched_noshuffle [1]}),
    .mi({open_n24923,\picorv32_core/mem_16bit_buffer [1]}),
    .fx({open_n24928,\picorv32_core/mem_rdata_latched [1]}),
    .q({open_n24929,\picorv32_core/mem_rdata_q [1]}));  // ../src/picorv32.v(508)
  // ../src/picorv32.v(508)
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("A*~C*~B*~D+A*~C*B*~D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000010101010),
    .INIT_LUTF1(16'b0000000000001010),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b1111111111111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b10|picorv32_core/reg0_b11  (
    .a({\picorv32_core/mem_rdata_q [10],\picorv32_core/mem_rdata_q [11]}),
    .c({\picorv32_core/mem_xfer_placeOpt_2 ,_al_u1464_o}),
    .clk(clk_pad),
    .d({_al_u1560_o,_al_u1560_o}),
    .e({_al_u1444_o,\picorv32_core/mem_xfer_placeOpt_2 }),
    .q({\picorv32_core/mem_rdata_q [10],\picorv32_core/mem_rdata_q [11]}));  // ../src/picorv32.v(508)
  // ../src/picorv32.v(508)
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(~0*~(~A*~B*D)))"),
    //.LUTF1("~D*~A*~B*~C+D*~A*~B*~C+D*A*~B*~C+~D*~A*B*~C+D*~A*B*~C+~D*A*B*~C+D*A*B*~C+~D*~A*~B*C+D*~A*~B*C+D*A*~B*C+~D*~A*B*C+D*~A*B*C+~D*A*B*C+D*A*B*C"),
    //.LUTG0("~(~C*~(~1*~(~A*~B*D)))"),
    //.LUTG1("D*~A*~B*~C+D*A*~B*~C+D*~A*B*~C+D*A*B*~C+D*~A*~B*C+D*A*~B*C+D*~A*B*C+D*A*B*C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111011111111),
    .INIT_LUTF1(16'b1111111111011101),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b1111111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b14|picorv32_core/reg0_b30  (
    .a({_al_u2353_o,_al_u2360_o}),
    .b({_al_u2359_o,_al_u2359_o}),
    .c({open_n24953,_al_u2357_o}),
    .clk(clk_pad),
    .d({_al_u2462_o,_al_u2353_o}),
    .e({_al_u2457_o,_al_u2354_o}),
    .q({\picorv32_core/mem_rdata_q [14],\picorv32_core/mem_rdata_q [30]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0)*~((B*~C*D))+~A*0*~((B*~C*D))+~(~A)*0*(B*~C*D)+~A*0*(B*~C*D))"),
    //.LUT1("(~A*~(1)*~((B*~C*D))+~A*1*~((B*~C*D))+~(~A)*1*(B*~C*D)+~A*1*(B*~C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101010101),
    .INIT_LUT1(16'b0101110101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b15  (
    .a({_al_u1585_o,_al_u1585_o}),
    .b({_al_u1580_o,_al_u1580_o}),
    .c({_al_u1579_o,_al_u1579_o}),
    .clk(clk_pad),
    .d({_al_u1569_o,_al_u1569_o}),
    .mi({open_n24986,\picorv32_core/mem_rdata_latched [5]}),
    .q({open_n24993,\picorv32_core/mem_rdata_q [15]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0)*~((C*~D*B))+~A*0*~((C*~D*B))+~(~A)*0*(C*~D*B)+~A*0*(C*~D*B))"),
    //.LUT1("(~A*~(1)*~((C*~D*B))+~A*1*~((C*~D*B))+~(~A)*1*(C*~D*B)+~A*1*(C*~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b0101010111010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b17  (
    .a({_al_u1591_o,_al_u1591_o}),
    .b({_al_u1569_o,_al_u1569_o}),
    .c({_al_u1580_o,_al_u1580_o}),
    .clk(clk_pad),
    .d({_al_u1579_o,_al_u1579_o}),
    .mi({open_n25005,\picorv32_core/mem_rdata_latched [12]}),
    .q({open_n25012,\picorv32_core/mem_rdata_q [17]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~B*~(D)*~(A)+~B*D*~(A)+~(~B)*D*A+~B*D*A))*~(C)+~0*(~B*~(D)*~(A)+~B*D*~(A)+~(~B)*D*A+~B*D*A)*~(C)+~(~0)*(~B*~(D)*~(A)+~B*D*~(A)+~(~B)*D*A+~B*D*A)*C+~0*(~B*~(D)*~(A)+~B*D*~(A)+~(~B)*D*A+~B*D*A)*C)"),
    //.LUT1("~(~1*~((~B*~(D)*~(A)+~B*D*~(A)+~(~B)*D*A+~B*D*A))*~(C)+~1*(~B*~(D)*~(A)+~B*D*~(A)+~(~B)*D*A+~B*D*A)*~(C)+~(~1)*(~B*~(D)*~(A)+~B*D*~(A)+~(~B)*D*A+~B*D*A)*C+~1*(~B*~(D)*~(A)+~B*D*~(A)+~(~B)*D*A+~B*D*A)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000011100000),
    .INIT_LUT1(16'b0100111111101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b1_placeOpt_1  (
    .a({_al_u1088_o,_al_u1088_o}),
    .b({\picorv32_core/mem_rdata_latched_noshuffle [1],\picorv32_core/mem_rdata_latched_noshuffle [1]}),
    .c({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .ce(\picorv32_core/mem_xfer_placeOpt_3 ),
    .clk(clk_pad),
    .d({_al_u1276_o,_al_u1276_o}),
    .mi({open_n25023,\picorv32_core/mem_16bit_buffer [1]}),
    .fx({open_n25028,\picorv32_core/mem_rdata_latched$1$_placeOpt_1 }));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))*~(B)+~0*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*~(B)+~(~0)*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B+~0*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B)"),
    //.LUT1("~(~1*~((~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))*~(A)+~1*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*~(A)+~(~1)*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A+~1*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100110000001000),
    .INIT_LUT1(16'b0111111101011101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b1_placeOpt_2  (
    .a({\picorv32_core/mux4_b0_sel_is_0_o ,_al_u1088_o}),
    .b({_al_u1088_o,\picorv32_core/mux4_b0_sel_is_0_o }),
    .c({_al_u1276_o,_al_u1276_o}),
    .ce(\picorv32_core/mem_xfer_placeOpt_3 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched_noshuffle [1],\picorv32_core/mem_rdata_latched_noshuffle [1]}),
    .mi({open_n25041,\picorv32_core/mem_16bit_buffer [1]}),
    .fx({open_n25046,\picorv32_core/mem_rdata_latched$1$_placeOpt_2 }));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))*~(B)+~0*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*~(B)+~(~0)*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B+~0*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B)"),
    //.LUT1("~(~1*~((~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))*~(A)+~1*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*~(A)+~(~1)*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A+~1*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100110000001000),
    .INIT_LUT1(16'b0111111101011101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b1_placeOpt_3  (
    .a({\picorv32_core/mux4_b0_sel_is_0_o ,_al_u1088_o}),
    .b({_al_u1088_o,\picorv32_core/mux4_b0_sel_is_0_o }),
    .c({_al_u1276_o,_al_u1276_o}),
    .ce(\picorv32_core/mem_xfer_placeOpt_3 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched_noshuffle [1],\picorv32_core/mem_rdata_latched_noshuffle [1]}),
    .mi({open_n25059,\picorv32_core/mem_16bit_buffer [1]}),
    .fx({open_n25064,\picorv32_core/mem_rdata_latched$1$_placeOpt_3 }));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))*~(B)+~0*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*~(B)+~(~0)*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B+~0*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B)"),
    //.LUT1("~(~1*~((~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))*~(A)+~1*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*~(A)+~(~1)*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A+~1*(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100110000001000),
    .INIT_LUT1(16'b0111111101011101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b1_placeOpt_4  (
    .a({\picorv32_core/mux4_b0_sel_is_0_o ,_al_u1088_o}),
    .b({_al_u1088_o,\picorv32_core/mux4_b0_sel_is_0_o }),
    .c({_al_u1276_o,_al_u1276_o}),
    .ce(\picorv32_core/mem_xfer_placeOpt_3 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched_noshuffle [1],\picorv32_core/mem_rdata_latched_noshuffle [1]}),
    .mi({open_n25077,\picorv32_core/mem_16bit_buffer [1]}),
    .fx({open_n25082,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))*~(A)+~0*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)*~(A)+~(~0)*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)*A+~0*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)*A)"),
    //.LUT1("~(~1*~((~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))*~(A)+~1*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)*~(A)+~(~1)*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)*A+~1*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000010101000),
    .INIT_LUT1(16'b0111010111111101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b2  (
    .a({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .b({_al_u1088_o,_al_u1088_o}),
    .c({\picorv32_core/mem_rdata_latched_noshuffle [2],\picorv32_core/mem_rdata_latched_noshuffle [2]}),
    .ce(\picorv32_core/mem_xfer_placeOpt_4 ),
    .clk(clk_pad),
    .d({_al_u1270_o,_al_u1270_o}),
    .mi({open_n25095,\picorv32_core/mem_16bit_buffer [2]}),
    .fx({open_n25100,\picorv32_core/mem_rdata_latched [2]}),
    .q({open_n25101,\picorv32_core/mem_rdata_q [2]}));  // ../src/picorv32.v(508)
  // ../src/picorv32.v(508)
  // ../src/picorv32.v(508)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*~C*~A+~B*D*~C*~A+~B*D*C*~A+~B*~D*~C*A+~B*D*~C*A+~B*D*C*A"),
    //.LUTF1("~A*~D*~B*~C+~A*D*~B*~C+~A*~D*B*~C+~A*D*B*~C+~A*~D*~B*C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    //.LUTG0("~B*~D*~C*~A+B*~D*~C*~A+~B*D*~C*~A+B*D*~C*~A+~B*~D*C*~A+B*~D*C*~A+~B*D*C*~A+B*D*C*~A+~B*~D*~C*A+B*~D*~C*A+~B*D*~C*A+B*D*~C*A+~B*~D*C*A+B*~D*C*A+~B*D*C*A+B*D*C*A"),
    //.LUTG1("~A*D*~B*~C+~A*D*B*~C+~A*~D*~B*C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b1111010111110101),
    .INIT_LUTG0(16'b1111111111111111),
    .INIT_LUTG1(16'b1111010111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b20|picorv32_core/reg0_b21  (
    .a({_al_u2281_o,open_n25102}),
    .b({open_n25103,_al_u2268_o}),
    .c({_al_u2285_o,_al_u1569_o}),
    .clk(clk_pad),
    .d({_al_u2279_o,_al_u2279_o}),
    .e({_al_u1569_o,_al_u2276_o}),
    .q({\picorv32_core/mem_rdata_q [20],\picorv32_core/mem_rdata_q [21]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C)*~((A*~B))*~(D)*~(0)+C*~((A*~B))*~(D)*~(0)+~(C)*(A*~B)*~(D)*~(0)+C*(A*~B)*~(D)*~(0)+~(C)*~((A*~B))*D*~(0)+C*~((A*~B))*D*~(0)+C*(A*~B)*D*~(0)+~(C)*~((A*~B))*D*0+C*~((A*~B))*D*0)"),
    //.LUT1("(~(C)*~((A*~B))*~(D)*~(1)+C*~((A*~B))*~(D)*~(1)+~(C)*(A*~B)*~(D)*~(1)+C*(A*~B)*~(D)*~(1)+~(C)*~((A*~B))*D*~(1)+C*~((A*~B))*D*~(1)+C*(A*~B)*D*~(1)+~(C)*~((A*~B))*D*1+C*~((A*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110111111111),
    .INIT_LUT1(16'b1101110100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b22  (
    .a({_al_u2342_o,_al_u2342_o}),
    .b({_al_u2340_o,_al_u2340_o}),
    .c({_al_u2279_o,_al_u2279_o}),
    .clk(clk_pad),
    .d({_al_u1569_o,_al_u1569_o}),
    .mi({open_n25136,_al_u2337_o}),
    .q({open_n25143,\picorv32_core/mem_rdata_q [22]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(A*~(D*~(0*B))))"),
    //.LUT1("~(~C*~(A*~(D*~(1*B))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111010),
    .INIT_LUT1(16'b1111100011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b23  (
    .a({_al_u1569_o,_al_u1569_o}),
    .b({_al_u2334_o,_al_u2334_o}),
    .c({_al_u2335_o,_al_u2335_o}),
    .clk(clk_pad),
    .d({_al_u2333_o,_al_u2333_o}),
    .mi({open_n25155,_al_u1606_o}),
    .q({open_n25162,\picorv32_core/mem_rdata_q [23]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~(~A*C*~B*~D))"),
    //.LUT1("(~1*~(~A*C*~B*~D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111101111),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b25  (
    .a({_al_u2392_o,_al_u2392_o}),
    .b({_al_u2387_o,_al_u2387_o}),
    .c({_al_u2390_o,_al_u2390_o}),
    .clk(clk_pad),
    .d({_al_u2385_o,_al_u2385_o}),
    .mi({open_n25174,_al_u2393_o}),
    .q({open_n25181,\picorv32_core/mem_rdata_q [25]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D*~(A*~(~0*~B))))"),
    //.LUT1("~(~C*~(D*~(A*~(~1*~B))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011111110000),
    .INIT_LUT1(16'b1111010111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b28  (
    .a({_al_u2378_o,_al_u2378_o}),
    .b({_al_u2376_o,_al_u2376_o}),
    .c({_al_u2373_o,_al_u2373_o}),
    .clk(clk_pad),
    .d({_al_u2380_o,_al_u2380_o}),
    .mi({open_n25193,_al_u1481_o_placeOpt_1}),
    .q({open_n25200,\picorv32_core/mem_rdata_q [28]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A))*~(B)+~0*(~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A)*~(B)+~(~0)*(~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A)*B+~0*(~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A)*B)"),
    //.LUT1("~(~1*~((~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A))*~(B)+~1*(~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A)*~(B)+~(~1)*(~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A)*B+~1*(~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000011001000),
    .INIT_LUT1(16'b0111001111111011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b3  (
    .a({_al_u1088_o,_al_u1088_o}),
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .c({\picorv32_core/mem_rdata_latched_noshuffle [3],\picorv32_core/mem_rdata_latched_noshuffle [3]}),
    .ce(\picorv32_core/mem_xfer_placeOpt_5 ),
    .clk(clk_pad),
    .d({_al_u1266_o,_al_u1266_o}),
    .mi({open_n25211,\picorv32_core/mem_16bit_buffer [3]}),
    .fx({open_n25216,\picorv32_core/mem_rdata_latched [3]}),
    .q({open_n25217,\picorv32_core/mem_rdata_q [3]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))*~(B)+~0*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*~(B)+~(~0)*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B+~0*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B)"),
    //.LUT1("~(~1*~((~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))*~(B)+~1*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*~(B)+~(~1)*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B+~1*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100110000001000),
    .INIT_LUT1(16'b0111111100111011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b4  (
    .a({_al_u1088_o,_al_u1088_o}),
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .c({_al_u1264_o,_al_u1264_o}),
    .ce(\picorv32_core/mem_xfer_placeOpt_4 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched_noshuffle [4],\picorv32_core/mem_rdata_latched_noshuffle [4]}),
    .mi({open_n25228,\picorv32_core/mem_16bit_buffer [4]}),
    .fx({open_n25233,\picorv32_core/mem_rdata_latched [4]}),
    .q({open_n25234,\picorv32_core/mem_rdata_q [4]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))*~(B)+~0*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*~(B)+~(~0)*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B+~0*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B)"),
    //.LUT1("~(~1*~((~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))*~(B)+~1*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*~(B)+~(~1)*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B+~1*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100110000001000),
    .INIT_LUT1(16'b0111111100111011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b6  (
    .a({_al_u1088_o,_al_u1088_o}),
    .b({\picorv32_core/mux4_b0_sel_is_0_o ,\picorv32_core/mux4_b0_sel_is_0_o }),
    .c({_al_u1257_o,_al_u1257_o}),
    .ce(\picorv32_core/mem_xfer_placeOpt_4 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched_noshuffle [6],\picorv32_core/mem_rdata_latched_noshuffle [6]}),
    .mi({open_n25245,\picorv32_core/mem_16bit_buffer [6]}),
    .fx({open_n25250,\picorv32_core/mem_rdata_latched [6]}),
    .q({open_n25251,\picorv32_core/mem_rdata_q [6]}));  // ../src/picorv32.v(508)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D)*~(B)*~(C)*~((0*A))+D*~(B)*~(C)*~((0*A))+~(D)*B*~(C)*~((0*A))+~(D)*~(B)*~(C)*(0*A)+D*~(B)*~(C)*(0*A)+~(D)*B*~(C)*(0*A)+D*B*~(C)*(0*A)+D*~(B)*C*(0*A)+D*B*C*(0*A))"),
    //.LUT1("(~(D)*~(A)*~(C)*~((1*B))+D*~(A)*~(C)*~((1*B))+~(D)*A*~(C)*~((1*B))+~(D)*~(A)*~(C)*(1*B)+D*~(A)*~(C)*(1*B)+~(D)*A*~(C)*(1*B)+D*A*~(C)*(1*B)+D*~(A)*C*(1*B)+D*A*C*(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100001111),
    .INIT_LUT1(16'b1100110100001111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg0_b7  (
    .a({_al_u1559_o,_al_u1532_o}),
    .b({_al_u1532_o,_al_u1559_o}),
    .c({_al_u1573_o,_al_u1573_o}),
    .clk(clk_pad),
    .d({_al_u1569_o,_al_u1569_o}),
    .mi({open_n25263,\picorv32_core/mem_rdata_latched [12]}),
    .q({open_n25270,\picorv32_core/mem_rdata_q [7]}));  // ../src/picorv32.v(508)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~D*B*~C+~A*D*B*~C+~A*~D*B*C+~A*D*B*C"),
    //.LUTF1("~A*~B*C*~D+~A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~D*B*~C+~A*D*B*~C+~A*~D*~B*C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    //.LUTG1("~A*~B*C*~D+~A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010001000100),
    .INIT_LUTF1(16'b1101110001010000),
    .INIT_LUTG0(16'b1111010011110100),
    .INIT_LUTG1(16'b1101110001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b10|picorv32_core/reg11_b9  (
    .a({_al_u896_o,_al_u896_o}),
    .b({\picorv32_core/decoded_imm_uj [10],\picorv32_core/mem_rdata_q [29]}),
    .c({\picorv32_core/mem_rdata_q [30],\picorv32_core/decoded_imm_uj [9]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_jal ,open_n25271}),
    .e({open_n25272,\picorv32_core/instr_jal }),
    .q(\picorv32_core/decoded_imm [10:9]));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(0*C)*~(D*~B))"),
    //.LUT1("~(~A*~(1*C)*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1111101111111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b12  (
    .a({_al_u908_o,_al_u908_o}),
    .b({_al_u665_o,_al_u665_o}),
    .c({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [12],\picorv32_core/mem_rdata_q [12]}),
    .mi({open_n25303,\picorv32_core/decoded_imm_uj [12]}),
    .q({open_n25310,\picorv32_core/decoded_imm [12]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(0*C)*~(D*~B))"),
    //.LUT1("~(~B*~(1*C)*~(D*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1111110111111100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b13  (
    .a({_al_u665_o,_al_u908_o}),
    .b({_al_u908_o,_al_u665_o}),
    .c({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [13],\picorv32_core/mem_rdata_q [13]}),
    .mi({open_n25321,\picorv32_core/decoded_imm_uj [13]}),
    .q({open_n25328,\picorv32_core/decoded_imm [13]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(0*C)*~(D*~B))"),
    //.LUT1("~(~A*~(1*C)*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1111101111111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b14  (
    .a({_al_u908_o,_al_u908_o}),
    .b({_al_u665_o,_al_u665_o}),
    .c({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [14],\picorv32_core/mem_rdata_q [14]}),
    .mi({open_n25339,\picorv32_core/decoded_imm_uj [14]}),
    .q({open_n25346,\picorv32_core/decoded_imm [14]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(0*C)*~(D*~B))"),
    //.LUT1("~(~A*~(1*D)*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1111111110111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b15  (
    .a({_al_u908_o,_al_u908_o}),
    .b({_al_u665_o,_al_u665_o}),
    .c({\picorv32_core/mem_rdata_q [15],\picorv32_core/instr_jal }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_jal ,\picorv32_core/mem_rdata_q [15]}),
    .mi({open_n25357,\picorv32_core/decoded_imm_uj [15]}),
    .q({open_n25364,\picorv32_core/decoded_imm [15]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(0*C)*~(D*~B))"),
    //.LUT1("~(~A*~(1*C)*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1111101111111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b16  (
    .a({_al_u908_o,_al_u908_o}),
    .b({_al_u665_o,_al_u665_o}),
    .c({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [16],\picorv32_core/mem_rdata_q [16]}),
    .mi({open_n25375,\picorv32_core/decoded_imm_uj [16]}),
    .q({open_n25382,\picorv32_core/decoded_imm [16]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(0*C)*~(D*~B))"),
    //.LUT1("~(~A*~(1*C)*~(B*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1111101011111110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b17  (
    .a({_al_u908_o,_al_u908_o}),
    .b({\picorv32_core/mem_rdata_q [17],_al_u665_o}),
    .c({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({_al_u665_o,\picorv32_core/mem_rdata_q [17]}),
    .mi({open_n25393,\picorv32_core/decoded_imm_uj [17]}),
    .q({open_n25400,\picorv32_core/decoded_imm [17]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(0*C)*~(D*~B))"),
    //.LUT1("~(~B*~(1*C)*~(A*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1111110011111110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b18  (
    .a({\picorv32_core/mem_rdata_q [18],_al_u908_o}),
    .b({_al_u908_o,_al_u665_o}),
    .c({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({_al_u665_o,\picorv32_core/mem_rdata_q [18]}),
    .mi({open_n25411,\picorv32_core/decoded_imm_uj [18]}),
    .q({open_n25418,\picorv32_core/decoded_imm [18]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(0*C)*~(D*~B))"),
    //.LUT1("~(~B*~(1*C)*~(A*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1111110011111110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b19  (
    .a({\picorv32_core/mem_rdata_q [19],_al_u908_o}),
    .b({_al_u908_o,_al_u665_o}),
    .c({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({_al_u665_o,\picorv32_core/mem_rdata_q [19]}),
    .mi({open_n25429,\picorv32_core/decoded_imm_uj [19]}),
    .q({open_n25436,\picorv32_core/decoded_imm [19]}));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~(~C*~B))*~(0*A))"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+B*~A*~C*D+B*A*~C*D+B*~A*C*D+B*A*C*D"),
    //.LUTG0("(~(D*~(~C*~B))*~(1*A))"),
    //.LUTG1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001111111111),
    .INIT_LUTF1(16'b1100110011111111),
    .INIT_LUTG0(16'b0000000101010101),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b1|_al_u933  (
    .a({open_n25437,\picorv32_core/instr_jal }),
    .b({\picorv32_core/mem_rdata_q [21],\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .c({open_n25438,\picorv32_core/is_sb_sh_sw }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({_al_u933_o,\picorv32_core/mem_rdata_q [8]}),
    .e({_al_u803_o,\picorv32_core/decoded_imm_uj [1]}),
    .f({open_n25454,_al_u933_o}),
    .q({\picorv32_core/decoded_imm [1],open_n25458}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(C*~(B*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0000111111001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b20|picorv32_core/reg11_b31  (
    .b({\picorv32_core/mem_rdata_q [20],_al_u665_o}),
    .c({_al_u909_o,\picorv32_core/mem_rdata_q [31]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({_al_u665_o,_al_u909_o}),
    .q({\picorv32_core/decoded_imm [20],\picorv32_core/decoded_imm [31]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(A*~B))"),
    //.LUT1("~(B*~(C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001011111111),
    .INIT_LUT1(16'b0011001111110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b21|picorv32_core/reg11_b30  (
    .a({open_n25479,\picorv32_core/mem_rdata_q [30]}),
    .b({_al_u909_o,_al_u665_o}),
    .c({\picorv32_core/mem_rdata_q [21],open_n25480}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({_al_u665_o,_al_u909_o}),
    .q({\picorv32_core/decoded_imm [21],\picorv32_core/decoded_imm [30]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~D*~A*~B+C*~D*~A*~B+~C*D*~A*~B+C*D*~A*~B+~C*~D*A*~B+C*~D*A*~B+~C*D*A*~B+C*D*A*~B+~C*~D*A*B+C*~D*A*B+~C*D*A*B+C*D*A*B"),
    //.LUTF1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+A*~D*~C*B+A*D*~C*B+A*~D*C*B+A*D*C*B"),
    //.LUTG0("~C*~D*~A*~B+C*~D*~A*~B+~C*D*~A*~B+C*D*~A*~B+~C*~D*A*~B+C*~D*A*~B+~C*D*A*~B+C*D*A*~B"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101110111011),
    .INIT_LUTF1(16'b1011101110111011),
    .INIT_LUTG0(16'b0011001100110011),
    .INIT_LUTG1(16'b0011001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b22|picorv32_core/reg11_b29  (
    .a({\picorv32_core/mem_rdata_q [22],\picorv32_core/mem_rdata_q [29]}),
    .b({_al_u909_o,_al_u909_o}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .e({_al_u665_o,_al_u665_o}),
    .q({\picorv32_core/decoded_imm [22],\picorv32_core/decoded_imm [29]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTF1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG0("~A*~B*D*~C+A*~B*D*~C+~A*~B*D*C+A*~B*D*C"),
    //.LUTG1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b1100110011111111),
    .INIT_LUTG0(16'b0011001100000000),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b23|picorv32_core/reg11_b28  (
    .b({\picorv32_core/mem_rdata_q [23],_al_u665_o}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({_al_u909_o,\picorv32_core/mem_rdata_q [28]}),
    .e({_al_u665_o,_al_u909_o}),
    .q({\picorv32_core/decoded_imm [23],\picorv32_core/decoded_imm [28]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~A))"),
    //.LUT1("~(D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b24|picorv32_core/reg11_b27  (
    .a({open_n25547,_al_u665_o}),
    .b({_al_u665_o,open_n25548}),
    .c({\picorv32_core/mem_rdata_q [24],\picorv32_core/mem_rdata_q [27]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({_al_u909_o,_al_u909_o}),
    .q({\picorv32_core/decoded_imm [24],\picorv32_core/decoded_imm [27]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~(C*~B))"),
    //.LUT1("~(A*~(B*~C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111010101110101),
    .INIT_LUT1(16'b0101110101011101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b25|picorv32_core/reg11_b26  (
    .a({_al_u909_o,_al_u909_o}),
    .b({\picorv32_core/mem_rdata_q [25],_al_u665_o}),
    .c({_al_u665_o,\picorv32_core/mem_rdata_q [26]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .q({\picorv32_core/decoded_imm [25],\picorv32_core/decoded_imm [26]}));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~(~C*~B))*~(0*A))"),
    //.LUTF1("~A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("(~(D*~(~C*~B))*~(1*A))"),
    //.LUTG1("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+~A*C*B*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001111111111),
    .INIT_LUTF1(16'b1111010111110101),
    .INIT_LUTG0(16'b0000000101010101),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b4|_al_u902  (
    .a({_al_u902_o,\picorv32_core/instr_jal }),
    .b({open_n25587,\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu }),
    .c({\picorv32_core/mem_rdata_q [24],\picorv32_core/is_sb_sh_sw }),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({open_n25588,\picorv32_core/mem_rdata_q [11]}),
    .e({_al_u803_o,\picorv32_core/decoded_imm_uj [4]}),
    .f({open_n25604,_al_u902_o}),
    .q({\picorv32_core/decoded_imm [4],open_n25608}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*C*~A+~B*D*C*~A+~B*~D*C*A+~B*D*C*A"),
    //.LUTF1("~B*~C*~A*D+~B*C*~A*D+~B*~C*A*D+~B*C*A*D"),
    //.LUTG0("~B*~D*C*~A+~B*D*C*~A+~B*~D*~C*A+B*~D*~C*A+~B*D*~C*A+B*D*~C*A+~B*~D*C*A+B*~D*C*A+~B*D*C*A+B*D*C*A"),
    //.LUTG1("~B*~C*A*~D+B*~C*A*~D+~B*C*A*~D+B*C*A*~D+~B*~C*~A*D+~B*C*~A*D+~B*~C*A*D+B*~C*A*D+~B*C*A*D+B*C*A*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000000110000),
    .INIT_LUTF1(16'b0011001100000000),
    .INIT_LUTG0(16'b1011101010111010),
    .INIT_LUTG1(16'b1011101110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b5|picorv32_core/reg11_b8  (
    .a({\picorv32_core/decoded_imm_uj [5],\picorv32_core/decoded_imm_uj [8]}),
    .b({_al_u896_o,_al_u896_o}),
    .c({open_n25609,\picorv32_core/mem_rdata_q [28]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_q [25],open_n25610}),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .q({\picorv32_core/decoded_imm [5],\picorv32_core/decoded_imm [8]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*~A))"),
    //.LUT1("~(~(B*D)*~(A*~C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110001010000),
    .INIT_LUT1(16'b1100111000001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg11_b6|picorv32_core/reg11_b7  (
    .a({\picorv32_core/mem_rdata_q [26],_al_u896_o}),
    .b({\picorv32_core/decoded_imm_uj [6],\picorv32_core/instr_jal }),
    .c({_al_u896_o,\picorv32_core/mem_rdata_q [27]}),
    .ce(\picorv32_core/n274 ),
    .clk(clk_pad),
    .d({\picorv32_core/instr_jal ,\picorv32_core/decoded_imm_uj [7]}),
    .q({\picorv32_core/decoded_imm [6],\picorv32_core/decoded_imm [7]}));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(B*~(C*(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100110011001100),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000110010001100),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg12_b1|_al_u1330  (
    .a({_al_u1330_o,\picorv32_core/n523_lutinv }),
    .b({open_n25649,_al_u1329_o}),
    .c({open_n25650,\picorv32_core/n664_lutinv_placeOpt_6 }),
    .clk(clk_pad),
    .d({open_n25652,\picorv32_core/cpuregs_rs2 [1]}),
    .e({resetn_placeOpt_17,\picorv32_core/decoded_rs2 [1]}),
    .f({open_n25668,_al_u1330_o}),
    .q({\picorv32_core/reg_sh [1],open_n25672}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(B*~A)"),
    //.LUTG0("(B*~(C*(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100110011001100),
    .INIT_LUTF1(16'b0100010001000100),
    .INIT_LUTG0(16'b0000110010001100),
    .INIT_LUTG1(16'b0100010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg12_b2|_al_u1325  (
    .a({_al_u1325_o,\picorv32_core/n523_lutinv }),
    .b({resetn_placeOpt_17,_al_u1324_o}),
    .c({open_n25673,\picorv32_core/n664_lutinv_placeOpt_6 }),
    .clk(clk_pad),
    .d({open_n25675,\picorv32_core/cpuregs_rs2 [2]}),
    .e({open_n25676,\picorv32_core/decoded_rs2 [2]}),
    .f({open_n25692,_al_u1325_o}),
    .q({\picorv32_core/reg_sh [2],open_n25696}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b0  (
    .a({\picorv32_core/n669_lutinv ,\picorv32_core/n669_lutinv }),
    .b({_al_u1904_o,_al_u1904_o}),
    .c({_al_u1900_o,_al_u1900_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25708,resetn_placeOpt_10}),
    .q({open_n25715,\picorv32_core/reg_out [0]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b11  (
    .a({\picorv32_core/n669_lutinv ,\picorv32_core/n669_lutinv }),
    .b({_al_u1881_o,_al_u1881_o}),
    .c({_al_u1877_o,_al_u1877_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25727,resetn_placeOpt_10}),
    .q({open_n25734,\picorv32_core/reg_out [11]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b12  (
    .a({\picorv32_core/n669_lutinv_placeOpt_1 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .b({_al_u1874_o,_al_u1874_o}),
    .c({_al_u1870_o,_al_u1870_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25746,resetn_placeOpt_12}),
    .q({open_n25753,\picorv32_core/reg_out [12]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*C*D)))"),
    //.LUT1("(1*~(B*~(A*C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1011001100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b15  (
    .a({\picorv32_core/n669_lutinv_placeOpt_1 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .b({_al_u1853_o,_al_u1853_o}),
    .c({_al_u1849_o,_al_u1849_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25765,resetn_placeOpt_12}),
    .q({open_n25772,\picorv32_core/reg_out [15]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b16  (
    .a({\picorv32_core/n669_lutinv ,\picorv32_core/n669_lutinv }),
    .b({_al_u1846_o,_al_u1846_o}),
    .c({_al_u1842_o,_al_u1842_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25784,resetn_placeOpt_10}),
    .q({open_n25791,\picorv32_core/reg_out [16]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b19  (
    .a({\picorv32_core/n669_lutinv ,\picorv32_core/n669_lutinv }),
    .b({_al_u1825_o,_al_u1825_o}),
    .c({_al_u1821_o,_al_u1821_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25803,resetn_placeOpt_10}),
    .q({open_n25810,\picorv32_core/reg_out [19]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b2  (
    .a({\picorv32_core/n669_lutinv ,\picorv32_core/n669_lutinv }),
    .b({_al_u1818_o,_al_u1818_o}),
    .c({_al_u1814_o,_al_u1814_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25822,resetn_placeOpt_10}),
    .q({open_n25829,\picorv32_core/reg_out [2]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b22  (
    .a({\picorv32_core/n669_lutinv_placeOpt_1 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .b({_al_u1794_o,_al_u1794_o}),
    .c({_al_u1790_o,_al_u1790_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25841,resetn_placeOpt_13}),
    .q({open_n25848,\picorv32_core/reg_out [22]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b23  (
    .a({\picorv32_core/n669_lutinv_placeOpt_1 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .b({_al_u1787_o,_al_u1787_o}),
    .c({_al_u1783_o,_al_u1783_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25860,resetn_placeOpt_12}),
    .q({open_n25867,\picorv32_core/reg_out [23]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b26  (
    .a({\picorv32_core/n669_lutinv_placeOpt_1 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .b({_al_u1766_o,_al_u1766_o}),
    .c({_al_u1762_o,_al_u1762_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25879,resetn_placeOpt_12}),
    .q({open_n25886,\picorv32_core/reg_out [26]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b27  (
    .a({\picorv32_core/n669_lutinv_placeOpt_1 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .b({_al_u1759_o,_al_u1759_o}),
    .c({_al_u1755_o,_al_u1755_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25898,resetn_placeOpt_12}),
    .q({open_n25905,\picorv32_core/reg_out [27]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b3  (
    .a({\picorv32_core/n669_lutinv ,\picorv32_core/n669_lutinv }),
    .b({_al_u1738_o,_al_u1738_o}),
    .c({_al_u1734_o,_al_u1734_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25917,resetn_placeOpt_10}),
    .q({open_n25924,\picorv32_core/reg_out [3]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b30  (
    .a({\picorv32_core/n669_lutinv_placeOpt_1 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .b({_al_u1727_o,_al_u1727_o}),
    .c({_al_u1723_o,_al_u1723_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25936,resetn_placeOpt_12}),
    .q({open_n25943,\picorv32_core/reg_out [30]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b5  (
    .a({\picorv32_core/n669_lutinv ,\picorv32_core/n669_lutinv }),
    .b({_al_u1701_o,_al_u1701_o}),
    .c({_al_u1697_o,_al_u1697_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25955,resetn_placeOpt_13}),
    .q({open_n25962,\picorv32_core/reg_out [5]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b6  (
    .a({\picorv32_core/n669_lutinv_placeOpt_1 ,\picorv32_core/n669_lutinv_placeOpt_1 }),
    .b({_al_u1692_o,_al_u1692_o}),
    .c({_al_u1688_o,_al_u1688_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25974,resetn_placeOpt_13}),
    .q({open_n25981,\picorv32_core/reg_out [6]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(B*~(A*~C*D)))"),
    //.LUT1("(1*~(B*~(A*~C*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0011101100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg13_b9  (
    .a({\picorv32_core/n669_lutinv ,\picorv32_core/n669_lutinv }),
    .b({_al_u1669_o,_al_u1669_o}),
    .c({_al_u1665_o,_al_u1665_o}),
    .clk(clk_pad),
    .d({\picorv32_core/n580 ,\picorv32_core/n580 }),
    .mi({open_n25993,resetn_placeOpt_10}),
    .q({open_n26000,\picorv32_core/reg_out [9]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b10  (
    .a({\picorv32_core/n434 [10],\picorv32_core/n434 [10]}),
    .b({\picorv32_core/n433 [10],\picorv32_core/n433 [10]}),
    .c({_al_u831_o,_al_u831_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26012,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26019,\picorv32_core/alu_out_q [10]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b11  (
    .a({\picorv32_core/n434 [11],\picorv32_core/n434 [11]}),
    .b({\picorv32_core/n433 [11],\picorv32_core/n433 [11]}),
    .c({_al_u833_o,_al_u833_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26031,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26038,\picorv32_core/alu_out_q [11]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b14  (
    .a({\picorv32_core/n434 [14],\picorv32_core/n434 [14]}),
    .b({\picorv32_core/n433 [14],\picorv32_core/n433 [14]}),
    .c({_al_u839_o,_al_u839_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26050,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26057,\picorv32_core/alu_out_q [14]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b15  (
    .a({\picorv32_core/n434 [15],\picorv32_core/n434 [15]}),
    .b({\picorv32_core/n433 [15],\picorv32_core/n433 [15]}),
    .c({_al_u841_o,_al_u841_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26069,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26076,\picorv32_core/alu_out_q [15]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b18  (
    .a({\picorv32_core/n434 [18],\picorv32_core/n434 [18]}),
    .b({\picorv32_core/n433 [18],\picorv32_core/n433 [18]}),
    .c({_al_u847_o,_al_u847_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26088,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26095,\picorv32_core/alu_out_q [18]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b19  (
    .a({\picorv32_core/n434 [19],\picorv32_core/n434 [19]}),
    .b({\picorv32_core/n433 [19],\picorv32_core/n433 [19]}),
    .c({_al_u849_o,_al_u849_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26107,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26114,\picorv32_core/alu_out_q [19]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b21  (
    .a({\picorv32_core/n434 [21],\picorv32_core/n434 [21]}),
    .b({\picorv32_core/n433 [21],\picorv32_core/n433 [21]}),
    .c({_al_u855_o,_al_u855_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26126,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26133,\picorv32_core/alu_out_q [21]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b22  (
    .a({\picorv32_core/n434 [22],\picorv32_core/n434 [22]}),
    .b({\picorv32_core/n433 [22],\picorv32_core/n433 [22]}),
    .c({_al_u857_o,_al_u857_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26145,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26152,\picorv32_core/alu_out_q [22]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b25  (
    .a({\picorv32_core/n434 [25],\picorv32_core/n434 [25]}),
    .b({\picorv32_core/n433 [25],\picorv32_core/n433 [25]}),
    .c({_al_u863_o,_al_u863_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26164,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26171,\picorv32_core/alu_out_q [25]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b26  (
    .a({\picorv32_core/n434 [26],\picorv32_core/n434 [26]}),
    .b({\picorv32_core/n433 [26],\picorv32_core/n433 [26]}),
    .c({_al_u865_o,_al_u865_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26183,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26190,\picorv32_core/alu_out_q [26]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b29  (
    .a({\picorv32_core/n434 [29],\picorv32_core/n434 [29]}),
    .b({\picorv32_core/n433 [29],\picorv32_core/n433 [29]}),
    .c({_al_u871_o,_al_u871_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26202,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26209,\picorv32_core/alu_out_q [29]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b3  (
    .a({\picorv32_core/n434 [3],\picorv32_core/n434 [3]}),
    .b({\picorv32_core/n433 [3],\picorv32_core/n433 [3]}),
    .c({_al_u873_o,_al_u873_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26221,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26228,\picorv32_core/alu_out_q [3]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b4  (
    .a({\picorv32_core/n434 [4],\picorv32_core/n434 [4]}),
    .b({\picorv32_core/n433 [4],\picorv32_core/n433 [4]}),
    .c({_al_u879_o,_al_u879_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26240,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26247,\picorv32_core/alu_out_q [4]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b5  (
    .a({\picorv32_core/n434 [5],\picorv32_core/n434 [5]}),
    .b({\picorv32_core/n433 [5],\picorv32_core/n433 [5]}),
    .c({_al_u881_o,_al_u881_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26259,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26266,\picorv32_core/alu_out_q [5]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b8  (
    .a({\picorv32_core/n434 [8],\picorv32_core/n434 [8]}),
    .b({\picorv32_core/n433 [8],\picorv32_core/n433 [8]}),
    .c({_al_u887_o,_al_u887_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26278,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26285,\picorv32_core/alu_out_q [8]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("~(~C*~(1*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111110011111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg14_b9  (
    .a({\picorv32_core/n434 [9],\picorv32_core/n434 [9]}),
    .b({\picorv32_core/n433 [9],\picorv32_core/n433 [9]}),
    .c({_al_u889_o,_al_u889_o}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_sub ,\picorv32_core/instr_sub }),
    .mi({open_n26297,\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub }),
    .q({open_n26304,\picorv32_core/alu_out_q [9]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+~A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+~A*~B*D*C+~A*B*D*C"),
    //.LUTF1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+~A*D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+~A*D*C*B"),
    //.LUTG0("~A*~B*~D*~C+A*~B*~D*~C+~A*~B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*~B*D*C"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+~A*D*C*~B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010111111111),
    .INIT_LUTF1(16'b0101111101011111),
    .INIT_LUTG0(16'b0001000100110011),
    .INIT_LUTG1(16'b0001001100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b11|picorv32_core/reg15_b8  (
    .a({\picorv32_core/instr_rdcycle ,\picorv32_core/instr_rdcycle }),
    .b({\picorv32_core/count_instr [43],\picorv32_core/instr_rdinstrh }),
    .c({\picorv32_core/count_cycle [11],open_n26305}),
    .clk(clk_pad),
    .d({open_n26307,\picorv32_core/count_cycle [8]}),
    .e({\picorv32_core/instr_rdinstrh ,\picorv32_core/count_instr [40]}),
    .mi({\picorv32_core/n459 [11],\picorv32_core/n459 [8]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1878_o,_al_u1674_o}),
    .q({\picorv32_core/count_cycle [11],\picorv32_core/count_cycle [8]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101111101011111),
    .INIT_LUTF1(16'b0011001111111111),
    .INIT_LUTG0(16'b0001001100010011),
    .INIT_LUTG1(16'b0001000101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b12|picorv32_core/reg15_b6  (
    .a({\picorv32_core/instr_rdcycle ,\picorv32_core/instr_rdcycle }),
    .b({\picorv32_core/instr_rdinstrh ,\picorv32_core/instr_rdinstrh }),
    .c({open_n26323,\picorv32_core/count_cycle [6]}),
    .clk(clk_pad),
    .d({\picorv32_core/count_instr [44],open_n26325}),
    .e({\picorv32_core/count_cycle [12],\picorv32_core/count_instr [38]}),
    .mi({\picorv32_core/n459 [12],\picorv32_core/n459 [6]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1871_o,_al_u1690_o}),
    .q({\picorv32_core/count_cycle [12],\picorv32_core/count_cycle [6]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b15|picorv32_core/reg15_b5  (
    .a({\picorv32_core/instr_rdcycle ,\picorv32_core/instr_rdcycle }),
    .b({\picorv32_core/count_cycle [15],\picorv32_core/instr_rdinstrh }),
    .c({\picorv32_core/instr_rdinstrh ,\picorv32_core/count_cycle [5]}),
    .clk(clk_pad),
    .d({\picorv32_core/count_instr [47],\picorv32_core/count_instr [37]}),
    .mi({\picorv32_core/n459 [15],\picorv32_core/n459 [5]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1850_o,_al_u1698_o}),
    .q({\picorv32_core/count_cycle [15],\picorv32_core/count_cycle [5]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b17|picorv32_core/reg15_b48  (
    .a({\picorv32_core/instr_rdcycle ,\picorv32_core/instr_rdcycleh }),
    .b({\picorv32_core/count_cycle [17],\picorv32_core/instr_rdinstr }),
    .c({\picorv32_core/instr_rdinstrh ,\picorv32_core/count_cycle [48]}),
    .clk(clk_pad),
    .d({\picorv32_core/count_instr [49],\picorv32_core/count_instr [16]}),
    .mi({\picorv32_core/n459 [17],\picorv32_core/n459 [48]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1836_o,_al_u1843_o}),
    .q({\picorv32_core/count_cycle [17],\picorv32_core/count_cycle [48]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+C*B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*~B*A*D+C*~B*A*D"),
    //.LUTF1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*~B*D*C+A*~B*D*C"),
    //.LUTG0("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+C*B*~A*~D+~C*~B*~A*D+C*~B*~A*D"),
    //.LUTG1("~A*~B*~D*~C+~A*B*~D*~C+~A*~B*D*~C+~A*B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111111111),
    .INIT_LUTF1(16'b0011111100111111),
    .INIT_LUTG0(16'b0001000101010101),
    .INIT_LUTG1(16'b0001010100010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b21|picorv32_core/reg15_b3  (
    .a({\picorv32_core/instr_rdcycle ,\picorv32_core/count_cycle [3]}),
    .b({\picorv32_core/instr_rdinstrh ,\picorv32_core/instr_rdinstrh }),
    .c({\picorv32_core/count_instr [53],open_n26369}),
    .clk(clk_pad),
    .d({open_n26371,\picorv32_core/count_instr [35]}),
    .e({\picorv32_core/count_cycle [21],\picorv32_core/instr_rdcycle }),
    .mi({\picorv32_core/n459 [21],\picorv32_core/n459 [3]}),
    .sr(resetn_placeOpt_5),
    .f({_al_u1798_o,_al_u1735_o}),
    .q({\picorv32_core/count_cycle [21],\picorv32_core/count_cycle [3]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+~A*B*~D*C+~A*~B*D*C+~A*B*D*C"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*~D*~C+A*~B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101111101011111),
    .INIT_LUTF1(16'b0101010111111111),
    .INIT_LUTG0(16'b0001001100010011),
    .INIT_LUTG1(16'b0001000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b22|picorv32_core/reg15_b29  (
    .a({\picorv32_core/instr_rdinstrh ,\picorv32_core/instr_rdinstrh }),
    .b({\picorv32_core/instr_rdcycle ,\picorv32_core/instr_rdcycle }),
    .c({open_n26387,\picorv32_core/count_instr [61]}),
    .clk(clk_pad),
    .d({\picorv32_core/count_instr [54],open_n26389}),
    .e({\picorv32_core/count_cycle [22],\picorv32_core/count_cycle [29]}),
    .mi({\picorv32_core/n459 [22],\picorv32_core/n459 [29]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1791_o,_al_u1743_o}),
    .q({\picorv32_core/count_cycle [22],\picorv32_core/count_cycle [29]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b23|picorv32_core/reg15_b27  (
    .a({\picorv32_core/instr_rdcycle ,\picorv32_core/instr_rdcycle }),
    .b({\picorv32_core/count_cycle [23],\picorv32_core/instr_rdinstrh }),
    .c({\picorv32_core/instr_rdinstrh ,\picorv32_core/count_cycle [27]}),
    .clk(clk_pad),
    .d({\picorv32_core/count_instr [55],\picorv32_core/count_instr [59]}),
    .mi({\picorv32_core/n459 [23],\picorv32_core/n459 [27]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1784_o,_al_u1756_o}),
    .q({\picorv32_core/count_cycle [23],\picorv32_core/count_cycle [27]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(B*D)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b24|picorv32_core/reg15_b25  (
    .a({\picorv32_core/instr_rdcycle ,\picorv32_core/instr_rdcycle }),
    .b({\picorv32_core/count_instr [56],\picorv32_core/instr_rdinstrh }),
    .c({\picorv32_core/count_cycle [24],\picorv32_core/count_cycle [25]}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_rdinstrh ,\picorv32_core/count_instr [57]}),
    .mi({\picorv32_core/n459 [24],\picorv32_core/n459 [25]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1777_o,_al_u1770_o}),
    .q({\picorv32_core/count_cycle [24],\picorv32_core/count_cycle [25]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(A*B)*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b33|picorv32_core/reg15_b63  (
    .a({\picorv32_core/count_instr [1],\picorv32_core/instr_rdcycleh }),
    .b({\picorv32_core/instr_rdinstr ,\picorv32_core/instr_rdinstr }),
    .c({\picorv32_core/count_cycle [33],\picorv32_core/count_cycle [63]}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_rdcycleh ,\picorv32_core/count_instr [31]}),
    .mi({\picorv32_core/n459 [33],\picorv32_core/n459 [63]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1892_o,_al_u1718_o}),
    .q({\picorv32_core/count_cycle [33],\picorv32_core/count_cycle [63]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(A*B)*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b36|picorv32_core/reg15_b62  (
    .a({\picorv32_core/count_instr [4],\picorv32_core/instr_rdcycleh }),
    .b({\picorv32_core/instr_rdinstr ,\picorv32_core/instr_rdinstr }),
    .c({\picorv32_core/count_cycle [36],\picorv32_core/count_cycle [62]}),
    .clk(clk_pad),
    .d({\picorv32_core/instr_rdcycleh ,\picorv32_core/count_instr [30]}),
    .mi({\picorv32_core/n459 [36],\picorv32_core/n459 [62]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1707_o,_al_u1725_o}),
    .q({\picorv32_core/count_cycle [36],\picorv32_core/count_cycle [62]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~D*~B+A*~C*~D*~B+~A*C*~D*~B+A*C*~D*~B+~A*~C*D*~B+~A*C*D*~B+~A*~C*~D*B+A*~C*~D*B+~A*C*~D*B+A*C*~D*B+~A*~C*D*B+~A*C*D*B"),
    //.LUTF1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG0("~A*~C*~D*~B+A*~C*~D*~B+~A*C*~D*~B+A*C*~D*~B+~A*~C*D*~B+~A*C*D*~B"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010111111111),
    .INIT_LUTF1(16'b0111011101110111),
    .INIT_LUTG0(16'b0001000100110011),
    .INIT_LUTG1(16'b0000000001110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b39|picorv32_core/reg15_b60  (
    .a({\picorv32_core/instr_rdcycleh ,\picorv32_core/instr_rdcycleh }),
    .b({\picorv32_core/count_cycle [39],\picorv32_core/count_instr [28]}),
    .clk(clk_pad),
    .d({\picorv32_core/count_instr [7],\picorv32_core/count_cycle [60]}),
    .e({\picorv32_core/instr_rdinstr ,\picorv32_core/instr_rdinstr }),
    .mi({\picorv32_core/n459 [39],\picorv32_core/n459 [60]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1680_o,_al_u1750_o}),
    .q({\picorv32_core/count_cycle [39],\picorv32_core/count_cycle [60]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b41|picorv32_core/reg15_b58  (
    .a({\picorv32_core/instr_rdcycleh ,\picorv32_core/instr_rdcycleh }),
    .b({\picorv32_core/instr_rdinstr ,\picorv32_core/instr_rdinstr }),
    .c({\picorv32_core/count_cycle [41],\picorv32_core/count_cycle [58]}),
    .clk(clk_pad),
    .d({\picorv32_core/count_instr [9],\picorv32_core/count_instr [26]}),
    .mi({\picorv32_core/n459 [41],\picorv32_core/n459 [58]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1666_o,_al_u1763_o}),
    .q({\picorv32_core/count_cycle [41],\picorv32_core/count_cycle [58]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b42|picorv32_core/reg15_b52  (
    .a({\picorv32_core/instr_rdcycleh ,\picorv32_core/instr_rdcycleh }),
    .b({\picorv32_core/instr_rdinstr ,\picorv32_core/instr_rdinstr }),
    .c({\picorv32_core/count_cycle [42],\picorv32_core/count_cycle [52]}),
    .clk(clk_pad),
    .d({\picorv32_core/count_instr [10],\picorv32_core/count_instr [20]}),
    .mi({\picorv32_core/n459 [42],\picorv32_core/n459 [52]}),
    .sr(resetn_placeOpt_14),
    .f({_al_u1885_o,_al_u1805_o}),
    .q({\picorv32_core/count_cycle [42],\picorv32_core/count_cycle [52]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTF1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*~B*D*C+A*~B*D*C"),
    //.LUTG0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG1("~A*~B*~D*~C+~A*B*~D*~C+~A*~B*D*~C+~A*B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111111111),
    .INIT_LUTF1(16'b0011111100111111),
    .INIT_LUTG0(16'b0001000101010101),
    .INIT_LUTG1(16'b0001010100010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b45|picorv32_core/reg15_b51  (
    .a({\picorv32_core/instr_rdcycleh ,\picorv32_core/instr_rdcycleh }),
    .b({\picorv32_core/instr_rdinstr ,\picorv32_core/instr_rdinstr }),
    .c({\picorv32_core/count_instr [13],open_n26507}),
    .clk(clk_pad),
    .d({open_n26509,\picorv32_core/count_instr [19]}),
    .e({\picorv32_core/count_cycle [45],\picorv32_core/count_cycle [51]}),
    .mi({\picorv32_core/n459 [45],\picorv32_core/n459 [51]}),
    .sr(resetn_placeOpt_4),
    .f({_al_u1864_o,_al_u1822_o}),
    .q({\picorv32_core/count_cycle [45],\picorv32_core/count_cycle [51]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~A*~C*~B+D*~A*~C*~B+~D*A*~C*~B+D*A*~C*~B+~D*~A*C*~B+D*~A*C*~B+~D*A*C*~B+D*A*C*~B+~D*~A*~C*B+D*~A*~C*B+~D*~A*C*B+D*~A*C*B"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*~A*~C*D+B*~A*~C*D+~B*~A*C*D+B*~A*C*D"),
    //.LUTG0("~D*~A*~C*~B+D*~A*~C*~B+~D*A*~C*~B+D*A*~C*~B+~D*~A*~C*B+D*~A*~C*B"),
    //.LUTG1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*~C*D+B*~A*~C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011101110111),
    .INIT_LUTF1(16'b0101010111111111),
    .INIT_LUTG0(16'b0000011100000111),
    .INIT_LUTG1(16'b0000010100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg15_b46|picorv32_core/reg15_b50  (
    .a({\picorv32_core/instr_rdinstr ,\picorv32_core/instr_rdinstr }),
    .b({open_n26525,\picorv32_core/count_instr [18]}),
    .c({\picorv32_core/count_cycle [46],\picorv32_core/count_cycle [50]}),
    .clk(clk_pad),
    .d({\picorv32_core/count_instr [14],open_n26527}),
    .e({\picorv32_core/instr_rdcycleh ,\picorv32_core/instr_rdcycleh }),
    .mi({\picorv32_core/n459 [46],\picorv32_core/n459 [50]}),
    .sr(resetn_placeOpt_4),
    .f({_al_u1857_o,_al_u1829_o}),
    .q({\picorv32_core/count_cycle [46],\picorv32_core/count_cycle [50]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D"),
    //.LUTF1("(B*~((A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0))*~(D)+B*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*~(D)+~(B)*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*D+B*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*D)"),
    //.LUTG0("A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("(B*~((A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1))*~(D)+B*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*~(D)+~(B)*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*D+B*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111010100100000),
    .INIT_LUTF1(16'b1010101011001100),
    .INIT_LUTG0(16'b1111110110101000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b0|picorv32_core/reg17_b0  (
    .a({\picorv32_core/n502 [0],\picorv32_core/sel15_b0_sel_is_3_o }),
    .b({\picorv32_core/n500 [0],\picorv32_core/latched_stalu }),
    .c({\picorv32_core/n504 [0],\picorv32_core/reg_out [0]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoder_trigger ,\picorv32_core/reg_next_pc [0]}),
    .e({\picorv32_core/instr_jal ,\picorv32_core/alu_out_q [0]}),
    .sr(resetn_placeOpt_7),
    .f({open_n26557,\picorv32_core/n500 [0]}),
    .q({\picorv32_core/reg_next_pc [0],\picorv32_core/reg_pc [0]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(A*~((B*~(D)*~(0)+B*D*~(0)+~(B)*D*0+B*D*0))*~(C)+A*(B*~(D)*~(0)+B*D*~(0)+~(B)*D*0+B*D*0)*~(C)+~(A)*(B*~(D)*~(0)+B*D*~(0)+~(B)*D*0+B*D*0)*C+A*(B*~(D)*~(0)+B*D*~(0)+~(B)*D*0+B*D*0)*C)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(A*~((B*~(D)*~(1)+B*D*~(1)+~(B)*D*1+B*D*1))*~(C)+A*(B*~(D)*~(1)+B*D*~(1)+~(B)*D*1+B*D*1)*~(C)+~(A)*(B*~(D)*~(1)+B*D*~(1)+~(B)*D*1+B*D*1)*C+A*(B*~(D)*~(1)+B*D*~(1)+~(B)*D*1+B*D*1)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1100101011001010),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b10|picorv32_core/reg18_b8  (
    .a({\picorv32_core/n500 [10],\picorv32_core/n502 [8]}),
    .b({\picorv32_core/n502 [10],\picorv32_core/n504 [8]}),
    .c({\picorv32_core/decoder_trigger ,\picorv32_core/n500 [8]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/n504 [10],\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [10],\picorv32_core/reg_next_pc [8]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(B*~((A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0))*~(D)+B*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*~(D)+~(B)*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*D+B*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*D)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(B*~((A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1))*~(D)+B*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*~(D)+~(B)*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*D+B*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1010101011001100),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b11|picorv32_core/reg18_b7  (
    .a({\picorv32_core/n502 [11],\picorv32_core/n502 [7]}),
    .b({\picorv32_core/n500 [11],\picorv32_core/n504 [7]}),
    .c({\picorv32_core/n504 [11],\picorv32_core/n500 [7]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoder_trigger ,\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [11],\picorv32_core/reg_next_pc [7]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(A*~((C*~(B)*~(0)+C*B*~(0)+~(C)*B*0+C*B*0))*~(D)+A*(C*~(B)*~(0)+C*B*~(0)+~(C)*B*0+C*B*0)*~(D)+~(A)*(C*~(B)*~(0)+C*B*~(0)+~(C)*B*0+C*B*0)*D+A*(C*~(B)*~(0)+C*B*~(0)+~(C)*B*0+C*B*0)*D)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(A*~((C*~(B)*~(1)+C*B*~(1)+~(C)*B*1+C*B*1))*~(D)+A*(C*~(B)*~(1)+C*B*~(1)+~(C)*B*1+C*B*1)*~(D)+~(A)*(C*~(B)*~(1)+C*B*~(1)+~(C)*B*1+C*B*1)*D+A*(C*~(B)*~(1)+C*B*~(1)+~(C)*B*1+C*B*1)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1111000010101010),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1100110010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b12|picorv32_core/reg18_b6  (
    .a({\picorv32_core/n500 [12],\picorv32_core/n502 [6]}),
    .b({\picorv32_core/n504 [12],\picorv32_core/n504 [6]}),
    .c({\picorv32_core/n502 [12],\picorv32_core/n500 [6]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoder_trigger ,\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [12],\picorv32_core/reg_next_pc [6]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(B*~((A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0))*~(D)+B*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*~(D)+~(B)*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*D+B*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*D)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(B*~((A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1))*~(D)+B*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*~(D)+~(B)*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*D+B*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1010101011001100),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b13|picorv32_core/reg18_b5  (
    .a({\picorv32_core/n502 [13],\picorv32_core/n502 [5]}),
    .b({\picorv32_core/n500 [13],\picorv32_core/n504 [5]}),
    .c({\picorv32_core/n504 [13],\picorv32_core/n500 [5]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoder_trigger ,\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [13],\picorv32_core/reg_next_pc [5]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(B*~((A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0))*~(C)+B*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*~(C)+~(B)*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*C+B*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*C)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(B*~((A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1))*~(C)+B*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*~(C)+~(B)*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*C+B*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1010110010101100),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b14|picorv32_core/reg18_b4  (
    .a({\picorv32_core/n502 [14],\picorv32_core/n502 [4]}),
    .b({\picorv32_core/n500 [14],\picorv32_core/n504 [4]}),
    .c({\picorv32_core/decoder_trigger ,\picorv32_core/n500 [4]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/n504 [14],\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [14],\picorv32_core/reg_next_pc [4]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(A*~((C*~(B)*~(0)+C*B*~(0)+~(C)*B*0+C*B*0))*~(D)+A*(C*~(B)*~(0)+C*B*~(0)+~(C)*B*0+C*B*0)*~(D)+~(A)*(C*~(B)*~(0)+C*B*~(0)+~(C)*B*0+C*B*0)*D+A*(C*~(B)*~(0)+C*B*~(0)+~(C)*B*0+C*B*0)*D)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(A*~((C*~(B)*~(1)+C*B*~(1)+~(C)*B*1+C*B*1))*~(D)+A*(C*~(B)*~(1)+C*B*~(1)+~(C)*B*1+C*B*1)*~(D)+~(A)*(C*~(B)*~(1)+C*B*~(1)+~(C)*B*1+C*B*1)*D+A*(C*~(B)*~(1)+C*B*~(1)+~(C)*B*1+C*B*1)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1111000010101010),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1100110010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b15|picorv32_core/reg18_b31  (
    .a({\picorv32_core/n500 [15],\picorv32_core/n502 [31]}),
    .b({\picorv32_core/n504 [15],\picorv32_core/n504 [31]}),
    .c({\picorv32_core/n502 [15],\picorv32_core/n500 [31]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoder_trigger ,\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [15],\picorv32_core/reg_next_pc [31]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(B*~((A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0))*~(D)+B*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*~(D)+~(B)*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*D+B*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*D)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(B*~((A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1))*~(D)+B*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*~(D)+~(B)*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*D+B*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1010101011001100),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b16|picorv32_core/reg18_b30  (
    .a({\picorv32_core/n502 [16],\picorv32_core/n502 [30]}),
    .b({\picorv32_core/n500 [16],\picorv32_core/n504 [30]}),
    .c({\picorv32_core/n504 [16],\picorv32_core/n500 [30]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoder_trigger ,\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [16],\picorv32_core/reg_next_pc [30]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(B*~((A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0))*~(C)+B*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*~(C)+~(B)*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*C+B*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*C)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(B*~((A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1))*~(C)+B*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*~(C)+~(B)*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*C+B*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1010110010101100),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b17|picorv32_core/reg18_b3  (
    .a({\picorv32_core/n502 [17],\picorv32_core/n502 [3]}),
    .b({\picorv32_core/n500 [17],\picorv32_core/n504 [3]}),
    .c({\picorv32_core/decoder_trigger ,\picorv32_core/n500 [3]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/n504 [17],\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [17],\picorv32_core/reg_next_pc [3]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(B*~((A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0))*~(D)+B*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*~(D)+~(B)*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*D+B*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*D)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(B*~((A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1))*~(D)+B*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*~(D)+~(B)*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*D+B*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1010101011001100),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b18|picorv32_core/reg18_b29  (
    .a({\picorv32_core/n502 [18],\picorv32_core/n502 [29]}),
    .b({\picorv32_core/n500 [18],\picorv32_core/n504 [29]}),
    .c({\picorv32_core/n504 [18],\picorv32_core/n500 [29]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoder_trigger ,\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [18],\picorv32_core/reg_next_pc [29]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(A*~((B*~(D)*~(0)+B*D*~(0)+~(B)*D*0+B*D*0))*~(C)+A*(B*~(D)*~(0)+B*D*~(0)+~(B)*D*0+B*D*0)*~(C)+~(A)*(B*~(D)*~(0)+B*D*~(0)+~(B)*D*0+B*D*0)*C+A*(B*~(D)*~(0)+B*D*~(0)+~(B)*D*0+B*D*0)*C)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(A*~((B*~(D)*~(1)+B*D*~(1)+~(B)*D*1+B*D*1))*~(C)+A*(B*~(D)*~(1)+B*D*~(1)+~(B)*D*1+B*D*1)*~(C)+~(A)*(B*~(D)*~(1)+B*D*~(1)+~(B)*D*1+B*D*1)*C+A*(B*~(D)*~(1)+B*D*~(1)+~(B)*D*1+B*D*1)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1100101011001010),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b19|picorv32_core/reg18_b28  (
    .a({\picorv32_core/n500 [19],\picorv32_core/n502 [28]}),
    .b({\picorv32_core/n502 [19],\picorv32_core/n504 [28]}),
    .c({\picorv32_core/decoder_trigger ,\picorv32_core/n500 [28]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/n504 [19],\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [19],\picorv32_core/reg_next_pc [28]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(B*~((A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0))*~(C)+B*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*~(C)+~(B)*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*C+B*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*C)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(B*~((A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1))*~(C)+B*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*~(C)+~(B)*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*C+B*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1010110010101100),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b1|picorv32_core/reg18_b27  (
    .a({\picorv32_core/n502 [1],\picorv32_core/n502 [27]}),
    .b({\picorv32_core/n500 [1],\picorv32_core/n504 [27]}),
    .c({\picorv32_core/decoder_trigger ,\picorv32_core/n500 [27]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/n504 [1],\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [1],\picorv32_core/reg_next_pc [27]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(B*~((A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0))*~(C)+B*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*~(C)+~(B)*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*C+B*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*C)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(B*~((A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1))*~(C)+B*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*~(C)+~(B)*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*C+B*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1010110010101100),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b20|picorv32_core/reg18_b26  (
    .a({\picorv32_core/n502 [20],\picorv32_core/n502 [26]}),
    .b({\picorv32_core/n500 [20],\picorv32_core/n504 [26]}),
    .c({\picorv32_core/decoder_trigger ,\picorv32_core/n500 [26]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/n504 [20],\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [20],\picorv32_core/reg_next_pc [26]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(A*~((B*~(D)*~(0)+B*D*~(0)+~(B)*D*0+B*D*0))*~(C)+A*(B*~(D)*~(0)+B*D*~(0)+~(B)*D*0+B*D*0)*~(C)+~(A)*(B*~(D)*~(0)+B*D*~(0)+~(B)*D*0+B*D*0)*C+A*(B*~(D)*~(0)+B*D*~(0)+~(B)*D*0+B*D*0)*C)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(A*~((B*~(D)*~(1)+B*D*~(1)+~(B)*D*1+B*D*1))*~(C)+A*(B*~(D)*~(1)+B*D*~(1)+~(B)*D*1+B*D*1)*~(C)+~(A)*(B*~(D)*~(1)+B*D*~(1)+~(B)*D*1+B*D*1)*C+A*(B*~(D)*~(1)+B*D*~(1)+~(B)*D*1+B*D*1)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1100101011001010),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b21|picorv32_core/reg18_b25  (
    .a({\picorv32_core/n500 [21],\picorv32_core/n502 [25]}),
    .b({\picorv32_core/n502 [21],\picorv32_core/n504 [25]}),
    .c({\picorv32_core/decoder_trigger ,\picorv32_core/n500 [25]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/n504 [21],\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [21],\picorv32_core/reg_next_pc [25]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(B*~((A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0))*~(C)+B*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*~(C)+~(B)*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*C+B*(A*~(D)*~(0)+A*D*~(0)+~(A)*D*0+A*D*0)*C)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(B*~((A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1))*~(C)+B*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*~(C)+~(B)*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*C+B*(A*~(D)*~(1)+A*D*~(1)+~(A)*D*1+A*D*1)*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1010110010101100),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b22|picorv32_core/reg18_b24  (
    .a({\picorv32_core/n502 [22],\picorv32_core/n502 [24]}),
    .b({\picorv32_core/n500 [22],\picorv32_core/n504 [24]}),
    .c({\picorv32_core/decoder_trigger ,\picorv32_core/n500 [24]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/n504 [22],\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [22],\picorv32_core/reg_next_pc [24]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0))*~(D)+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*~(D)+~(C)*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D+C*(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)*D)"),
    //.LUTF1("(B*~((A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0))*~(D)+B*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*~(D)+~(B)*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*D+B*(A*~(C)*~(0)+A*C*~(0)+~(A)*C*0+A*C*0)*D)"),
    //.LUTG0("(C*~((A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1))*~(D)+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*~(D)+~(C)*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D+C*(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)*D)"),
    //.LUTG1("(B*~((A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1))*~(D)+B*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*~(D)+~(B)*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*D+B*(A*~(C)*~(1)+A*C*~(1)+~(A)*C*1+A*C*1)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b1010101011001100),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("SET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg18_b2|picorv32_core/reg18_b23  (
    .a({\picorv32_core/n502 [2],\picorv32_core/n502 [23]}),
    .b({\picorv32_core/n500 [2],\picorv32_core/n504 [23]}),
    .c({\picorv32_core/n504 [2],\picorv32_core/n500 [23]}),
    .ce(\picorv32_core/n663 ),
    .clk(clk_pad),
    .d({\picorv32_core/decoder_trigger ,\picorv32_core/decoder_trigger }),
    .e({\picorv32_core/instr_jal ,\picorv32_core/instr_jal }),
    .sr(resetn_placeOpt_7),
    .q({\picorv32_core/reg_next_pc [2],\picorv32_core/reg_next_pc [23]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b10|picorv32_core/reg19_b9  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi(\picorv32_core/n503 [10:9]),
    .sr(resetn_placeOpt_5),
    .q(\picorv32_core/count_instr [10:9]));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b11|picorv32_core/reg19_b8  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [11],\picorv32_core/n503 [8]}),
    .sr(resetn_placeOpt_5),
    .q({\picorv32_core/count_instr [11],\picorv32_core/count_instr [8]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b12|picorv32_core/reg19_b7  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [12],\picorv32_core/n503 [7]}),
    .sr(resetn_placeOpt_5),
    .q({\picorv32_core/count_instr [12],\picorv32_core/count_instr [7]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b13|picorv32_core/reg19_b63  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [13],\picorv32_core/n503 [63]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [13],\picorv32_core/count_instr [63]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b14|picorv32_core/reg19_b62  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [14],\picorv32_core/n503 [62]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [14],\picorv32_core/count_instr [62]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b15|picorv32_core/reg19_b61  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [15],\picorv32_core/n503 [61]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [15],\picorv32_core/count_instr [61]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b16|picorv32_core/reg19_b60  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [16],\picorv32_core/n503 [60]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [16],\picorv32_core/count_instr [60]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b17|picorv32_core/reg19_b6  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [17],\picorv32_core/n503 [6]}),
    .sr(resetn_placeOpt_5),
    .q({\picorv32_core/count_instr [17],\picorv32_core/count_instr [6]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b18|picorv32_core/reg19_b59  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [18],\picorv32_core/n503 [59]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [18],\picorv32_core/count_instr [59]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b19|picorv32_core/reg19_b58  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [19],\picorv32_core/n503 [58]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [19],\picorv32_core/count_instr [58]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b20|picorv32_core/reg19_b57  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [20],\picorv32_core/n503 [57]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [20],\picorv32_core/count_instr [57]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b21|picorv32_core/reg19_b56  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [21],\picorv32_core/n503 [56]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [21],\picorv32_core/count_instr [56]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b22|picorv32_core/reg19_b55  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [22],\picorv32_core/n503 [55]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [22],\picorv32_core/count_instr [55]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b23|picorv32_core/reg19_b54  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [23],\picorv32_core/n503 [54]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [23],\picorv32_core/count_instr [54]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b24|picorv32_core/reg19_b53  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [24],\picorv32_core/n503 [53]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [24],\picorv32_core/count_instr [53]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b25|picorv32_core/reg19_b52  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [25],\picorv32_core/n503 [52]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [25],\picorv32_core/count_instr [52]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b26|picorv32_core/reg19_b51  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [26],\picorv32_core/n503 [51]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [26],\picorv32_core/count_instr [51]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b27|picorv32_core/reg19_b50  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [27],\picorv32_core/n503 [50]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [27],\picorv32_core/count_instr [50]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b28|picorv32_core/reg19_b5  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [28],\picorv32_core/n503 [5]}),
    .sr(resetn_placeOpt_5),
    .q({\picorv32_core/count_instr [28],\picorv32_core/count_instr [5]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b29|picorv32_core/reg19_b49  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [29],\picorv32_core/n503 [49]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [29],\picorv32_core/count_instr [49]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b2|picorv32_core/reg19_b48  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [2],\picorv32_core/n503 [48]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [2],\picorv32_core/count_instr [48]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b30|picorv32_core/reg19_b47  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [30],\picorv32_core/n503 [47]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [30],\picorv32_core/count_instr [47]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b31|picorv32_core/reg19_b46  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [31],\picorv32_core/n503 [46]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [31],\picorv32_core/count_instr [46]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b34|picorv32_core/reg19_b45  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [34],\picorv32_core/n503 [45]}),
    .sr(resetn_placeOpt_14),
    .q({\picorv32_core/count_instr [34],\picorv32_core/count_instr [45]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b35|picorv32_core/reg19_b44  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [35],\picorv32_core/n503 [44]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [35],\picorv32_core/count_instr [44]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b36|picorv32_core/reg19_b43  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [36],\picorv32_core/n503 [43]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [36],\picorv32_core/count_instr [43]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b37|picorv32_core/reg19_b42  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [37],\picorv32_core/n503 [42]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [37],\picorv32_core/count_instr [42]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b38|picorv32_core/reg19_b41  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [38],\picorv32_core/n503 [41]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [38],\picorv32_core/count_instr [41]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b39|picorv32_core/reg19_b40  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [39],\picorv32_core/n503 [40]}),
    .sr(resetn_placeOpt_4),
    .q({\picorv32_core/count_instr [39],\picorv32_core/count_instr [40]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \picorv32_core/reg19_b3|picorv32_core/reg19_b4  (
    .ce(\picorv32_core/sel39_b0_sel_is_3_o ),
    .clk(clk_pad),
    .mi({\picorv32_core/n503 [3],\picorv32_core/n503 [4]}),
    .sr(resetn_placeOpt_5),
    .q({\picorv32_core/count_instr [3],\picorv32_core/count_instr [4]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C*~(~0*B*~D)))"),
    //.LUT1("(A*~(C*~(~1*B*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101010001010),
    .INIT_LUT1(16'b0000101000001010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg1_b1  (
    .a({_al_u1615_o,_al_u1615_o}),
    .b({_al_u1577_o,_al_u1577_o}),
    .c({_al_u1614_o,_al_u1614_o}),
    .clk(clk_pad),
    .d({\picorv32_core/mem_la_read ,\picorv32_core/mem_la_read }),
    .mi({open_n27607,\picorv32_core/mem_do_rinst }),
    .q({open_n27614,\picorv32_core/mem_state [1]}));  // ../src/picorv32.v(605)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*A*~C+~D*B*A*~C+~D*~B*A*C+~D*B*A*C"),
    //.LUTF1("~A*C*~B*~D+A*C*~B*~D+~A*C*B*~D+A*C*B*~D"),
    //.LUTG0("~D*B*~A*~C+D*B*~A*~C+~D*~B*A*~C+~D*B*A*~C+D*B*A*~C+~D*B*~A*C+D*B*~A*C+~D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTG1("A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+A*~C*~B*D+A*C*~B*D+A*~C*B*D+A*C*B*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010101010),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1100110011101110),
    .INIT_LUTG1(16'b1010101011111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg24_b0|picorv32_core/reg24_b3  (
    .a({\picorv32_core/decoded_rd [0],\picorv32_core/latched_rd [3]}),
    .b({open_n27615,\picorv32_core/n663 }),
    .c({\picorv32_core/latched_rd [0],open_n27616}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1153_o,_al_u1153_o}),
    .e({\picorv32_core/n663 ,\picorv32_core/decoded_rd [3]}),
    .q({\picorv32_core/latched_rd [0],\picorv32_core/latched_rd [3]}));  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*~A))"),
    //.LUT1("~(~(C*B)*~(D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110001010000),
    .INIT_LUT1(16'b1101010111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg24_b1|picorv32_core/reg24_b2  (
    .a({_al_u1153_o,_al_u1153_o}),
    .b({\picorv32_core/n663 ,\picorv32_core/n663 }),
    .c({\picorv32_core/decoded_rd [1],\picorv32_core/latched_rd [2]}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/latched_rd [1],\picorv32_core/decoded_rd [2]}),
    .q({\picorv32_core/latched_rd [1],\picorv32_core/latched_rd [2]}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(D*~C)*~(B*~A))"),
    //.LUT1("~(1*~(D*~C)*~(B*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0100111101000100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b0  (
    .a({_al_u2258_o,_al_u2258_o}),
    .b({_al_u2259_o,_al_u2259_o}),
    .c({_al_u2260_o,_al_u2260_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2261_o,_al_u2261_o}),
    .mi({open_n27665,_al_u2265_o}),
    .q({open_n27672,\picorv32_core/pcpi_rs1$0$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(B*~A)*~(D*~C))"),
    //.LUT1("~(1*~(B*~A)*~(D*~C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0100111101000100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b10  (
    .a({_al_u2249_o,_al_u2249_o}),
    .b({_al_u2250_o,_al_u2250_o}),
    .c({_al_u2247_o,_al_u2247_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2248_o,_al_u2248_o}),
    .mi({open_n27683,_al_u2256_o}),
    .q({open_n27690,\picorv32_core/pcpi_rs1$10$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(B*~C)*~(D*~A))"),
    //.LUT1("~(1*~(B*~C)*~(D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0101110100001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b11  (
    .a({_al_u2236_o,_al_u2236_o}),
    .b({_al_u2239_o,_al_u2239_o}),
    .c({_al_u2238_o,_al_u2238_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2237_o,_al_u2237_o}),
    .mi({open_n27701,_al_u2245_o}),
    .q({open_n27708,\picorv32_core/pcpi_rs1$11$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(B*~A)*~(D*~C))"),
    //.LUT1("~(1*~(B*~A)*~(D*~C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0100111101000100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b14  (
    .a({_al_u2205_o,_al_u2205_o}),
    .b({_al_u2206_o,_al_u2206_o}),
    .c({_al_u2203_o,_al_u2203_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2204_o,_al_u2204_o}),
    .mi({open_n27719,_al_u2212_o}),
    .q({open_n27726,\picorv32_core/pcpi_rs1$14$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(C*~A)*~(B*~D))"),
    //.LUT1("~(1*~(C*~A)*~(B*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0101000011011100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b15  (
    .a({_al_u2194_o,_al_u2194_o}),
    .b({_al_u2193_o,_al_u2193_o}),
    .c({_al_u2195_o,_al_u2195_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2192_o,_al_u2192_o}),
    .mi({open_n27737,_al_u2201_o}),
    .q({open_n27744,\picorv32_core/pcpi_rs1$15$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(A*~B)*~(C*~D))"),
    //.LUT1("~(1*~(A*~B)*~(C*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0010001011110010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b18  (
    .a({_al_u2162_o,_al_u2162_o}),
    .b({_al_u2161_o,_al_u2161_o}),
    .c({_al_u2160_o,_al_u2160_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2159_o,_al_u2159_o}),
    .mi({open_n27755,_al_u2168_o}),
    .q({open_n27762,\picorv32_core/pcpi_rs1$18$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(B*~A)*~(D*~C))"),
    //.LUT1("~(1*~(B*~A)*~(D*~C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0100111101000100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b19  (
    .a({_al_u2150_o,_al_u2150_o}),
    .b({_al_u2151_o,_al_u2151_o}),
    .c({_al_u2148_o,_al_u2148_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2149_o,_al_u2149_o}),
    .mi({open_n27773,_al_u2157_o}),
    .q({open_n27780,\picorv32_core/pcpi_rs1$19$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(B*~A)*~(D*~C))"),
    //.LUT1("~(1*~(B*~A)*~(D*~C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0100111101000100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b2  (
    .a({_al_u2022_o,_al_u2022_o}),
    .b({_al_u2023_o,_al_u2023_o}),
    .c({_al_u2020_o,_al_u2020_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2021_o,_al_u2021_o}),
    .mi({open_n27791,_al_u2028_o}),
    .q({open_n27798,\picorv32_core/pcpi_rs1$2$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(C*~A)*~(B*~D))"),
    //.LUT1("~(1*~(C*~A)*~(B*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0101000011011100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b22  (
    .a({_al_u2107_o,_al_u2107_o}),
    .b({_al_u2106_o,_al_u2106_o}),
    .c({_al_u2108_o,_al_u2108_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2105_o,_al_u2105_o}),
    .mi({open_n27809,_al_u2114_o}),
    .q({open_n27816,\picorv32_core/pcpi_rs1$22$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(C*~A)*~(B*~D))"),
    //.LUT1("~(1*~(C*~A)*~(B*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0101000011011100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b23  (
    .a({_al_u2096_o,_al_u2096_o}),
    .b({_al_u2095_o,_al_u2095_o}),
    .c({_al_u2097_o,_al_u2097_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2094_o,_al_u2094_o}),
    .mi({open_n27827,_al_u2103_o}),
    .q({open_n27834,\picorv32_core/pcpi_rs1$23$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(C*~A)*~(B*~D))"),
    //.LUT1("~(1*~(C*~A)*~(B*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0101000011011100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b26  (
    .a({_al_u2063_o,_al_u2063_o}),
    .b({_al_u2062_o,_al_u2062_o}),
    .c({_al_u2064_o,_al_u2064_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2061_o,_al_u2061_o}),
    .mi({open_n27845,_al_u2070_o}),
    .q({open_n27852,\picorv32_core/pcpi_rs1$26$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(A*~C)*~(B*~D))"),
    //.LUT1("~(1*~(A*~C)*~(B*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0000101011001110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b27  (
    .a({_al_u2053_o,_al_u2053_o}),
    .b({_al_u2051_o,_al_u2051_o}),
    .c({_al_u2052_o,_al_u2052_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2050_o,_al_u2050_o}),
    .mi({open_n27863,_al_u2059_o}),
    .q({open_n27870,\picorv32_core/pcpi_rs1$27$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(C*~A)*~(B*~D))"),
    //.LUT1("~(1*~(C*~A)*~(B*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0101000011011100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b28  (
    .a({_al_u2042_o,_al_u2042_o}),
    .b({_al_u2041_o,_al_u2041_o}),
    .c({_al_u2043_o,_al_u2043_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2040_o,_al_u2040_o}),
    .mi({open_n27881,_al_u2048_o}),
    .q({open_n27888,\picorv32_core/pcpi_rs1$28$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(A*~C)*~(B*~D))"),
    //.LUT1("~(1*~(A*~C)*~(B*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0000101011001110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b3  (
    .a({_al_u1992_o,_al_u1992_o}),
    .b({_al_u1990_o,_al_u1990_o}),
    .c({_al_u1991_o,_al_u1991_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1989_o,_al_u1989_o}),
    .mi({open_n27899,_al_u1997_o}),
    .q({open_n27906,\picorv32_core/pcpi_rs1$3$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(D*~A)*~(B*~C))"),
    //.LUT1("~(1*~(D*~A)*~(B*~C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0101110100001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b31  (
    .a({_al_u2001_o,_al_u2001_o}),
    .b({_al_u2000_o,_al_u2000_o}),
    .c({_al_u1999_o,_al_u1999_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u2002_o,_al_u2002_o}),
    .mi({open_n27917,_al_u2007_o}),
    .q({open_n27924,\picorv32_core/pcpi_rs1$31$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(D*~B)*~(C*~A))"),
    //.LUT1("~(1*~(D*~B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0111001101010000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b5  (
    .a({_al_u1967_o,_al_u1967_o}),
    .b({_al_u1969_o,_al_u1969_o}),
    .c({_al_u1968_o,_al_u1968_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1970_o,_al_u1970_o}),
    .mi({open_n27935,_al_u1976_o}),
    .q({open_n27942,\picorv32_core/pcpi_rs1$5$ }));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("~(0*~(A*~C)*~(B*~D))"),
    //.LUT1("~(1*~(A*~C)*~(B*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111111),
    .INIT_LUT1(16'b0000101011001110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg25_b8  (
    .a({_al_u1937_o,_al_u1937_o}),
    .b({_al_u1935_o,_al_u1935_o}),
    .c({_al_u1936_o,_al_u1936_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1934_o,_al_u1934_o}),
    .mi({open_n27953,_al_u1943_o}),
    .q({open_n27960,\picorv32_core/pcpi_rs1$8$ }));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b1100110011111111),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b11|_al_u1423  (
    .a({open_n27961,\picorv32_core/n523_lutinv }),
    .b({\picorv32_core/cpuregs_rs2 [11],_al_u1339_o}),
    .c({open_n27962,\picorv32_core/n664_lutinv_placeOpt_2 }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1423_o,\picorv32_core/decoded_imm [11]}),
    .e({_al_u1337_o,\picorv32_core/pcpi_rs2$11$ }),
    .f({open_n27978,_al_u1423_o}),
    .q({\picorv32_core/pcpi_rs2$11$ ,open_n27982}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0000111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b12|_al_u1420  (
    .a({open_n27983,\picorv32_core/n523_lutinv }),
    .b({open_n27984,_al_u1339_o}),
    .c({_al_u1337_o,\picorv32_core/n664_lutinv }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1420_o,\picorv32_core/decoded_imm [12]}),
    .e({\picorv32_core/cpuregs_rs2 [12],\picorv32_core/pcpi_rs2$12$ }),
    .f({open_n28000,_al_u1420_o}),
    .q({\picorv32_core/pcpi_rs2$12$ ,open_n28004}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~(A*~(D*~B))"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~(A*~(D*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b0111011101010101),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b15|_al_u1411  (
    .a({_al_u1411_o,\picorv32_core/n523_lutinv }),
    .b({_al_u1337_o,_al_u1339_o}),
    .c({open_n28005,\picorv32_core/n664_lutinv }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_rs2 [15],\picorv32_core/decoded_imm [15]}),
    .e({open_n28006,\picorv32_core/pcpi_rs2$15$ }),
    .f({open_n28022,_al_u1411_o}),
    .q({\picorv32_core/pcpi_rs2$15$ ,open_n28026}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b1111010111110101),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b17|_al_u1405  (
    .a({_al_u1405_o,\picorv32_core/n523_lutinv }),
    .b({open_n28027,_al_u1339_o}),
    .c({\picorv32_core/cpuregs_rs2 [17],\picorv32_core/n664_lutinv }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({open_n28028,\picorv32_core/decoded_imm [17]}),
    .e({_al_u1337_o,\picorv32_core/pcpi_rs2$17$ }),
    .f({open_n28044,_al_u1405_o}),
    .q({\picorv32_core/pcpi_rs2$17$ ,open_n28048}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~(D*~(C*~A))"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~(D*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b0101000011111111),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0101000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b18|_al_u1402  (
    .a({_al_u1337_o,\picorv32_core/n523_lutinv }),
    .b({open_n28049,_al_u1339_o}),
    .c({\picorv32_core/cpuregs_rs2 [18],\picorv32_core/n664_lutinv }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1402_o,\picorv32_core/decoded_imm [18]}),
    .e({open_n28050,\picorv32_core/pcpi_rs2$18$ }),
    .f({open_n28066,_al_u1402_o}),
    .q({\picorv32_core/pcpi_rs2$18$ ,open_n28070}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*~B*C*A+D*~B*C*A"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b1011101110111011),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b0011001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b19|_al_u849  (
    .a({\picorv32_core/cpuregs_rs2 [19],_al_u826_o}),
    .b({_al_u1399_o,_al_u827_o}),
    .c({open_n28071,_al_u828_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({open_n28072,\picorv32_core/pcpi_rs1$19$ }),
    .e({_al_u1337_o,\picorv32_core/pcpi_rs2$19$ }),
    .f({open_n28088,_al_u849_o}),
    .q({\picorv32_core/pcpi_rs2$19$ ,open_n28092}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(B*(0*~(D)*~(C)+0*D*~(C)+~(0)*D*C+0*D*C)))"),
    //.LUTF1("D*~C*~A*~B+D*C*~A*~B+~D*~C*A*~B+D*~C*A*~B+~D*C*A*~B+D*C*A*~B+D*~C*~A*B+D*C*~A*B+~D*~C*A*B+D*~C*A*B+~D*C*A*B+D*C*A*B"),
    //.LUTG0("(~A*~(B*(1*~(D)*~(C)+1*D*~(C)+~(1)*D*C+1*D*C)))"),
    //.LUTG1("~D*~C*~A*~B+D*~C*~A*~B+D*C*~A*~B+~D*~C*A*~B+D*~C*A*~B+~D*C*A*~B+D*C*A*~B+~D*~C*~A*B+D*~C*~A*B+D*C*~A*B+~D*~C*A*B+D*~C*A*B+~D*C*A*B+D*C*A*B"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010101010101),
    .INIT_LUTF1(16'b1111111110101010),
    .INIT_LUTG0(16'b0001000101010001),
    .INIT_LUTG1(16'b1111111110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b1|_al_u1329  (
    .a({\picorv32_core/sel42_b1/B4 ,\picorv32_core/sel42_b1/B4 }),
    .b({open_n28093,\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv }),
    .c({_al_u1339_o,\picorv32_core/n554 }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/sel42_b1/B5 ,\picorv32_core/n559 [1]}),
    .e({mem_la_wdata[1],\picorv32_core/n564 [1]}),
    .f({open_n28109,_al_u1329_o}),
    .q({mem_la_wdata[1],open_n28113}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("~A*~B*~D*~C+A*~B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("~A*~B*~D*~C+A*~B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*~B*D*C+A*~B*D*C"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b1111111100110011),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b0011001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b21|_al_u855  (
    .a({open_n28114,_al_u826_o}),
    .b({_al_u1391_o,_al_u827_o}),
    .c({open_n28115,_al_u828_o}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_rs2 [21],\picorv32_core/pcpi_rs1$21$ }),
    .e({_al_u1337_o,\picorv32_core/pcpi_rs2$21$ }),
    .f({open_n28131,_al_u855_o}),
    .q({\picorv32_core/pcpi_rs2$21$ ,open_n28135}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~(D*~(A*~C))"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~(D*~(A*~C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b0000101011111111),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0000101011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b22|_al_u1388  (
    .a({\picorv32_core/cpuregs_rs2 [22],\picorv32_core/n523_lutinv }),
    .b({open_n28136,_al_u1339_o}),
    .c({_al_u1337_o,\picorv32_core/n664_lutinv_placeOpt_7 }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1388_o,\picorv32_core/decoded_imm [22]}),
    .e({open_n28137,\picorv32_core/pcpi_rs2$22$ }),
    .f({open_n28153,_al_u1388_o}),
    .q({\picorv32_core/pcpi_rs2$22$ ,open_n28157}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+~A*C*B*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b1101110111011101),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b23|_al_u1385  (
    .a({_al_u1385_o,\picorv32_core/n523_lutinv }),
    .b({\picorv32_core/cpuregs_rs2 [23],_al_u1339_o}),
    .c({open_n28158,\picorv32_core/n664_lutinv_placeOpt_3 }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({open_n28159,\picorv32_core/decoded_imm [23]}),
    .e({_al_u1337_o,\picorv32_core/pcpi_rs2$23$ }),
    .f({open_n28175,_al_u1385_o}),
    .q({\picorv32_core/pcpi_rs2$23$ ,open_n28179}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~(D*~(B*~A))"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~(D*~(B*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b0100010011111111),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0100010011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b26|_al_u1376  (
    .a({_al_u1337_o,\picorv32_core/n523_lutinv }),
    .b({\picorv32_core/cpuregs_rs2 [26],_al_u1339_o}),
    .c({open_n28180,\picorv32_core/n664_lutinv_placeOpt_4 }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1376_o,\picorv32_core/decoded_imm [26]}),
    .e({open_n28181,\picorv32_core/pcpi_rs2$26$ }),
    .f({open_n28197,_al_u1376_o}),
    .q({\picorv32_core/pcpi_rs2$26$ ,open_n28201}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b1111010111110101),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b27|_al_u1373  (
    .a({_al_u1373_o,\picorv32_core/n523_lutinv }),
    .b({open_n28202,_al_u1339_o}),
    .c({\picorv32_core/cpuregs_rs2 [27],\picorv32_core/n664_lutinv_placeOpt_7 }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({open_n28203,\picorv32_core/decoded_imm [27]}),
    .e({_al_u1337_o,\picorv32_core/pcpi_rs2$27$ }),
    .f({open_n28219,_al_u1373_o}),
    .q({\picorv32_core/pcpi_rs2$27$ ,open_n28223}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0101010111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b30|_al_u1362  (
    .a({_al_u1337_o,\picorv32_core/n523_lutinv }),
    .b({open_n28224,_al_u1339_o}),
    .c({open_n28225,\picorv32_core/n664_lutinv }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1362_o,\picorv32_core/decoded_imm [30]}),
    .e({\picorv32_core/cpuregs_rs2 [30],\picorv32_core/pcpi_rs2$30$ }),
    .f({open_n28241,_al_u1362_o}),
    .q({\picorv32_core/pcpi_rs2$30$ ,open_n28245}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*C*~B*D+A*C*~B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b1111000011111111),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b31|_al_u1359  (
    .a({open_n28246,\picorv32_core/n523_lutinv }),
    .b({open_n28247,_al_u1339_o}),
    .c({\picorv32_core/cpuregs_rs2 [31],\picorv32_core/n664_lutinv_placeOpt_7 }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1359_o,\picorv32_core/decoded_imm [31]}),
    .e({_al_u1337_o,\picorv32_core/pcpi_rs2$31$ }),
    .f({open_n28263,_al_u1359_o}),
    .q({\picorv32_core/pcpi_rs2$31$ ,open_n28267}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(B*(0*~(D)*~(C)+0*D*~(C)+~(0)*D*C+0*D*C)))"),
    //.LUTF1("A*~C*~B*~D+A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+A*~C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("(~A*~(B*(1*~(D)*~(C)+1*D*~(C)+~(1)*D*C+1*D*C)))"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+A*~C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010101010101),
    .INIT_LUTF1(16'b1110111011101110),
    .INIT_LUTG0(16'b0001000101010001),
    .INIT_LUTG1(16'b1110111011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b4|_al_u1315  (
    .a({\picorv32_core/sel42_b4/B5 ,\picorv32_core/sel42_b4/B4 }),
    .b({\picorv32_core/sel42_b4/B4 ,\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o_lutinv }),
    .c({open_n28268,\picorv32_core/n554 }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1339_o,\picorv32_core/n559 [4]}),
    .e({mem_la_wdata[4],\picorv32_core/n564 [4]}),
    .f({open_n28284,_al_u1315_o}),
    .q({mem_la_wdata[4],open_n28288}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b1111010111110101),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b5|_al_u1352  (
    .a({_al_u1352_o,\picorv32_core/n523_lutinv }),
    .b({open_n28289,_al_u1339_o}),
    .c({\picorv32_core/cpuregs_rs2 [5],\picorv32_core/n664_lutinv_placeOpt_7 }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({open_n28290,\picorv32_core/decoded_imm [5]}),
    .e({_al_u1337_o,mem_la_wdata[5]}),
    .f({open_n28306,_al_u1352_o}),
    .q({mem_la_wdata[5],open_n28310}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~(A*~(D*~B))"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~(A*~(D*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b0111011101010101),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b6|_al_u1349  (
    .a({_al_u1349_o,\picorv32_core/n523_lutinv }),
    .b({_al_u1337_o,_al_u1339_o}),
    .c({open_n28311,\picorv32_core/n664_lutinv_placeOpt_7 }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({\picorv32_core/cpuregs_rs2 [6],\picorv32_core/decoded_imm [6]}),
    .e({open_n28312,mem_la_wdata[6]}),
    .f({open_n28328,_al_u1349_o}),
    .q({mem_la_wdata[6],open_n28332}));  // ../src/picorv32.v(1906)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(0*~B)*~(D*C*~A))"),
    //.LUTF1("~(A*~(B*~D))"),
    //.LUTG0("(~(1*~B)*~(D*C*~A))"),
    //.LUTG1("~(A*~(B*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111111111111),
    .INIT_LUTF1(16'b0101010111011101),
    .INIT_LUTG0(16'b1000110011001100),
    .INIT_LUTG1(16'b0101010111011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg26_b8|_al_u1343  (
    .a({_al_u1343_o,\picorv32_core/n523_lutinv }),
    .b({\picorv32_core/cpuregs_rs2 [8],_al_u1339_o}),
    .c({open_n28333,\picorv32_core/n664_lutinv_placeOpt_2 }),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .d({_al_u1337_o,\picorv32_core/decoded_imm [8]}),
    .e({open_n28334,\picorv32_core/pcpi_rs2$8$ }),
    .f({open_n28350,_al_u1343_o}),
    .q({\picorv32_core/pcpi_rs2$8$ ,open_n28354}));  // ../src/picorv32.v(1906)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUT1("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010011000000),
    .INIT_LUT1(16'b1110111011001111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg5_b1  (
    .a({_al_u1089_o,_al_u1089_o}),
    .b({mem_rdata[17],mem_rdata[17]}),
    .c({\picorv32_core/mux51_b0_sel_is_3_o ,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_la_read ,\picorv32_core/mem_la_read }),
    .mi({open_n28365,\picorv32_core/mem_16bit_buffer [1]}),
    .q({open_n28372,\picorv32_core/mem_16bit_buffer [1]}));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUT1("(A*~(1)*~((~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C))+A*1*~((~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C))+~(A)*1*(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)+A*1*(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010011000000),
    .INIT_LUT1(16'b1110101011101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg5_b11  (
    .a({mem_rdata[27],_al_u1089_o}),
    .b({_al_u1089_o,mem_rdata[27]}),
    .c({\picorv32_core/mem_la_read ,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mux51_b0_sel_is_3_o ,\picorv32_core/mem_la_read }),
    .mi({open_n28383,\picorv32_core/mem_16bit_buffer [11]}),
    .q({open_n28390,\picorv32_core/mem_16bit_buffer [11]}));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUT1("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010011000000),
    .INIT_LUT1(16'b1110111011001111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg5_b12  (
    .a({_al_u1089_o,_al_u1089_o}),
    .b({mem_rdata[28],mem_rdata[28]}),
    .c({\picorv32_core/mux51_b0_sel_is_3_o ,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_la_read ,\picorv32_core/mem_la_read }),
    .mi({open_n28401,\picorv32_core/mem_16bit_buffer [12]}),
    .q({open_n28408,\picorv32_core/mem_16bit_buffer [12]}));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUT1("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010011000000),
    .INIT_LUT1(16'b1110111011001111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg5_b13  (
    .a({_al_u1089_o,_al_u1089_o}),
    .b({mem_rdata[29],mem_rdata[29]}),
    .c({\picorv32_core/mux51_b0_sel_is_3_o ,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_la_read ,\picorv32_core/mem_la_read }),
    .mi({open_n28419,\picorv32_core/mem_16bit_buffer [13]}),
    .q({open_n28426,\picorv32_core/mem_16bit_buffer [13]}));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUT1("(A*~(1)*~((~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D))+A*1*~((~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D))+~(A)*1*(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D)+A*1*(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010011000000),
    .INIT_LUT1(16'b1110111010101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg5_b14  (
    .a({mem_rdata[30],_al_u1089_o}),
    .b({_al_u1089_o,mem_rdata[30]}),
    .c({\picorv32_core/mux51_b0_sel_is_3_o ,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_la_read ,\picorv32_core/mem_la_read }),
    .mi({open_n28437,\picorv32_core/mem_16bit_buffer [14]}),
    .q({open_n28444,\picorv32_core/mem_16bit_buffer [14]}));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUT1("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010011000000),
    .INIT_LUT1(16'b1110111011001111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg5_b2  (
    .a({_al_u1089_o,_al_u1089_o}),
    .b({mem_rdata[18],mem_rdata[18]}),
    .c({\picorv32_core/mux51_b0_sel_is_3_o ,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_la_read ,\picorv32_core/mem_la_read }),
    .mi({open_n28455,\picorv32_core/mem_16bit_buffer [2]}),
    .q({open_n28462,\picorv32_core/mem_16bit_buffer [2]}));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUT1("(A*~(1)*~((~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C))+A*1*~((~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C))+~(A)*1*(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)+A*1*(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010011000000),
    .INIT_LUT1(16'b1110101011101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg5_b3  (
    .a({mem_rdata[19],_al_u1089_o}),
    .b({_al_u1089_o,mem_rdata[19]}),
    .c({\picorv32_core/mem_la_read ,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mux51_b0_sel_is_3_o ,\picorv32_core/mem_la_read }),
    .mi({open_n28473,\picorv32_core/mem_16bit_buffer [3]}),
    .q({open_n28480,\picorv32_core/mem_16bit_buffer [3]}));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUT1("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010011000000),
    .INIT_LUT1(16'b1110111011001111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg5_b5  (
    .a({_al_u1089_o,_al_u1089_o}),
    .b({mem_rdata[21],mem_rdata[21]}),
    .c({\picorv32_core/mux51_b0_sel_is_3_o ,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_la_read ,\picorv32_core/mem_la_read }),
    .mi({open_n28491,\picorv32_core/mem_16bit_buffer [5]}),
    .q({open_n28498,\picorv32_core/mem_16bit_buffer [5]}));  // ../src/picorv32.v(605)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*0*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*0*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUT1("(B*~(1)*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+B*1*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))+~(B)*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)+B*1*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010011000000),
    .INIT_LUT1(16'b1110111011001111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg5_b7  (
    .a({_al_u1089_o,_al_u1089_o}),
    .b({mem_rdata[23],mem_rdata[23]}),
    .c({\picorv32_core/mux51_b0_sel_is_3_o ,\picorv32_core/mux51_b0_sel_is_3_o }),
    .ce(\picorv32_core/mux68_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_la_read ,\picorv32_core/mem_la_read }),
    .mi({open_n28509,\picorv32_core/mem_16bit_buffer [7]}),
    .q({open_n28516,\picorv32_core/mem_16bit_buffer [7]}));  // ../src/picorv32.v(605)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A)*~((B*C))+D*A*~((B*C))+~(D)*A*(B*C)+D*A*(B*C))"),
    //.LUT1("(C*~(B)*~((A*D))+C*B*~((A*D))+~(C)*B*(A*D)+C*B*(A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111110000000),
    .INIT_LUT1(16'b1101100011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg6_b11|picorv32_core/reg6_b15  (
    .a({\picorv32_core/mem_rdata_latched [0],_al_u1481_o_placeOpt_4}),
    .b({\picorv32_core/mem_rdata_latched [20],\picorv32_core/mem_rdata_latched [0]}),
    .c({\picorv32_core/mem_rdata_latched [12],\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched$1$_placeOpt_4 ,\picorv32_core/mem_rdata_latched [12]}),
    .q({\picorv32_core/decoded_imm_uj [11],\picorv32_core/decoded_imm_uj [15]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("A*D*C*~B+A*D*C*B"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111100001110000),
    .INIT_LUTF1(16'b1010000000000000),
    .INIT_LUTG0(16'b1111100001110000),
    .INIT_LUTG1(16'b1111010111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg6_b14|picorv32_core/reg6_b13  (
    .a({\picorv32_core/mem_rdata_latched$0$_placeOpt_3 ,\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }),
    .b({open_n28535,\picorv32_core/mem_rdata_latched [1]}),
    .c({_al_u1483_o,\picorv32_core/mem_rdata_latched [12]}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched [1],_al_u1485_o}),
    .e({\picorv32_core/mem_rdata_latched [12],open_n28536}),
    .q(\picorv32_core/decoded_imm_uj [14:13]));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("C*~A*D*B+C*A*D*B"),
    //.LUTG0("~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG1("~C*~A*~D*~B+C*~A*~D*~B+~C*A*~D*~B+C*A*~D*~B+~C*~A*D*~B+C*~A*D*~B+~C*A*D*~B+C*A*D*~B+~C*~A*~D*B+~C*A*~D*B+~C*~A*D*B+C*~A*D*B+~C*A*D*B+C*A*D*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011001100),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1010110010101100),
    .INIT_LUTG1(16'b1111111100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg6_b3|picorv32_core/reg6_b6  (
    .a({open_n28557,\picorv32_core/mem_rdata_latched [26]}),
    .b({\picorv32_core/mem_rdata_latched$1$_placeOpt_4 ,\picorv32_core/mux79_b0/B0_3 }),
    .c({\picorv32_core/mem_rdata_latched$0$_placeOpt_3 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_rdata_latched [23],open_n28558}),
    .e({\picorv32_core/mem_rdata_latched [5],\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }),
    .q({\picorv32_core/decoded_imm_uj [3],\picorv32_core/decoded_imm_uj [6]}));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(~(B)*~(C)*~(D)*~(0)+B*~(C)*~(D)*~(0)+~(B)*C*~(D)*~(0)+B*C*~(D)*~(0)+~(B)*~(C)*D*~(0)+~(B)*C*D*~(0)+~(B)*C*~(D)*0+~(B)*C*D*0))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("(~A*(~(B)*~(C)*~(D)*~(1)+B*~(C)*~(D)*~(1)+~(B)*C*~(D)*~(1)+B*C*~(D)*~(1)+~(B)*~(C)*D*~(1)+~(B)*C*D*~(1)+~(B)*C*~(D)*1+~(B)*C*D*1))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001000101010101),
    .INIT_LUTF1(16'b0101010111011101),
    .INIT_LUTG0(16'b0001000000010000),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg7_b0|_al_u2294  (
    .a({_al_u2294_o,_al_u2292_o}),
    .b({_al_u1606_o,_al_u2293_o}),
    .c({open_n28579,\picorv32_core/n180 }),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u2290_o,\picorv32_core/mux81_sel_is_1_o }),
    .e({_al_u2297_o,\picorv32_core/mux79_b0/B0_3 }),
    .f({open_n28595,_al_u2294_o}),
    .q({\picorv32_core/decoded_rd [0],open_n28599}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(A*(~(C)*~(D)*~(B)*~(0)+C*~(D)*~(B)*~(0)+~(C)*D*~(B)*~(0)+C*D*~(B)*~(0)+~(C)*~(D)*B*~(0)+~(C)*D*B*~(0)+~(C)*~(D)*~(B)*0+C*~(D)*~(B)*0+~(C)*~(D)*B*0+C*~(D)*B*0+~(C)*D*B*0+C*D*B*0))"),
    //.LUT1("~(A*(~(C)*~(D)*~(B)*~(1)+C*~(D)*~(B)*~(1)+~(C)*D*~(B)*~(1)+C*D*~(B)*~(1)+~(C)*~(D)*B*~(1)+~(C)*D*B*~(1)+~(C)*~(D)*~(B)*1+C*~(D)*~(B)*1+~(C)*~(D)*B*1+C*~(D)*B*1+~(C)*D*B*1+C*D*B*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101010111010101),
    .INIT_LUT1(16'b0111011101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg7_b1  (
    .a({_al_u2455_o,_al_u2455_o}),
    .b({\picorv32_core/mem_rdata_latched [1],\picorv32_core/mem_rdata_latched [1]}),
    .c({_al_u2453_o,_al_u2453_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u2454_o,_al_u2454_o}),
    .mi({open_n28610,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .q({open_n28617,\picorv32_core/decoded_rd [1]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(A*(~(C)*~(D)*~(B)*~(0)+C*~(D)*~(B)*~(0)+~(C)*D*~(B)*~(0)+C*D*~(B)*~(0)+C*~(D)*B*~(0)+C*D*B*~(0)+~(C)*~(D)*~(B)*0+C*~(D)*~(B)*0+~(C)*~(D)*B*0+C*~(D)*B*0+~(C)*D*B*0+C*D*B*0))"),
    //.LUT1("~(A*(~(C)*~(D)*~(B)*~(1)+C*~(D)*~(B)*~(1)+~(C)*D*~(B)*~(1)+C*D*~(B)*~(1)+C*~(D)*B*~(1)+C*D*B*~(1)+~(C)*~(D)*~(B)*1+C*~(D)*~(B)*1+~(C)*~(D)*B*1+C*~(D)*B*1+~(C)*D*B*1+C*D*B*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101110101011101),
    .INIT_LUT1(16'b0111011101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg7_b2  (
    .a({_al_u2451_o,_al_u2451_o}),
    .b({\picorv32_core/mem_rdata_latched [1],\picorv32_core/mem_rdata_latched [1]}),
    .c({_al_u2449_o,_al_u2449_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u2450_o,_al_u2450_o}),
    .mi({open_n28628,\picorv32_core/mem_rdata_latched$0$_placeOpt_4 }),
    .q({open_n28635,\picorv32_core/decoded_rd [2]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~((~0*~(D)*~(B)+~0*D*~(B)+~(~0)*D*B+~0*D*B)*~(A*C))"),
    //.LUT1("~((~1*~(D)*~(A)+~1*D*~(A)+~(~1)*D*A+~1*D*A)*~(B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010000011101100),
    .INIT_LUT1(16'b1101010111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg8_b0  (
    .a({\picorv32_core/n180 ,\picorv32_core/mux79_b0/B0_3 }),
    .b({\picorv32_core/mux79_b0/B0_3 ,\picorv32_core/n180 }),
    .c({_al_u2427_o,_al_u2427_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u2441_o,_al_u2441_o}),
    .mi({open_n28646,_al_u1481_o_placeOpt_4}),
    .q({open_n28653,\picorv32_core/decoded_rs1 [0]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~((~0*~(D)*~(B)+~0*D*~(B)+~(~0)*D*B+~0*D*B)*~(A*C))"),
    //.LUT1("~((~1*~(D)*~(A)+~1*D*~(A)+~(~1)*D*A+~1*D*A)*~(B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010000011101100),
    .INIT_LUT1(16'b1101010111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg8_b2  (
    .a({\picorv32_core/n180 ,\picorv32_core/mux79_b2/B0_3 }),
    .b({\picorv32_core/mux79_b2/B0_3 ,\picorv32_core/n180 }),
    .c({_al_u2427_o,_al_u2427_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u2431_o,_al_u2431_o}),
    .mi({open_n28664,\picorv32_core/mem_rdata_latched [17]}),
    .q({open_n28671,\picorv32_core/decoded_rs1 [2]}));  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*~C*D+B*~A*~C*D+~B*A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTF1("C*~A*~B*~D+C*A*~B*~D+~C*~A*B*~D+C*~A*B*~D+~C*A*B*~D+C*A*B*~D+C*~A*~B*D+C*A*~B*D+~C*~A*B*D+C*~A*B*D+~C*A*B*D+C*A*B*D"),
    //.LUTG0("B*A*~C*~D+B*A*C*~D+~B*~A*~C*D+B*~A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+B*A*C*D"),
    //.LUTG1("~C*~A*~B*~D+C*~A*~B*~D+~C*A*~B*~D+C*A*~B*~D+~C*~A*B*~D+C*~A*B*~D+~C*A*B*~D+C*A*B*~D+~C*~A*B*D+C*~A*B*D+~C*A*B*D+C*A*B*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b1111110011111100),
    .INIT_LUTG0(16'b1101110110001000),
    .INIT_LUTG1(16'b1100110011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg8_b3|picorv32_core/reg6_b18  (
    .a({open_n28672,\picorv32_core/mem_rdata_latched [0]}),
    .b({_al_u2427_o,\picorv32_core/mem_rdata_latched [18]}),
    .c({\picorv32_core/mem_rdata_latched [18],open_n28673}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u2426_o,\picorv32_core/mem_rdata_latched [12]}),
    .e({\picorv32_core/n180 ,\picorv32_core/mem_rdata_latched$1$_placeOpt_4 }),
    .q({\picorv32_core/decoded_rs1 [3],\picorv32_core/decoded_imm_uj [18]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(0*~D*~(~A*~B)))"),
    //.LUT1("~(~D*~(1*~C*~(~A*~B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011110000),
    .INIT_LUT1(16'b1111111100001110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg8_b4  (
    .a({_al_u1606_o,_al_u1606_o}),
    .b({_al_u2293_o,_al_u2293_o}),
    .c({_al_u2420_o,_al_u2421_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u2421_o,_al_u2420_o}),
    .mi({open_n28704,_al_u2422_o}),
    .q({open_n28711,\picorv32_core/decoded_rs1 [4]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(~0*B*~(~A*~C)))"),
    //.LUT1("~(~D*~(~1*B*~(~A*~C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111001000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg9_b0  (
    .a({_al_u1627_o,_al_u1627_o}),
    .b({\picorv32_core/mem_rdata_latched [2],\picorv32_core/mem_rdata_latched [2]}),
    .c({_al_u1623_o,_al_u1623_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u1646_o,_al_u1646_o}),
    .mi({open_n28722,\picorv32_core/mem_rdata_latched [1]}),
    .q({open_n28729,\picorv32_core/decoded_rs2 [0]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(~0*A*~(~C*~D)))"),
    //.LUT1("~(~B*~(~1*A*~(~C*~D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111011101100),
    .INIT_LUT1(16'b1100110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg9_b1  (
    .a({\picorv32_core/mem_rdata_latched [3],\picorv32_core/mem_rdata_latched [3]}),
    .b({_al_u1643_o,_al_u1643_o}),
    .c({_al_u1627_o,_al_u1627_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u1623_o,_al_u1623_o}),
    .mi({open_n28740,\picorv32_core/mem_rdata_latched [1]}),
    .q({open_n28747,\picorv32_core/decoded_rs2 [1]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(~0*B*~(~A*~C)))"),
    //.LUT1("~(~D*~(~1*A*~(~B*~C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111001000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg9_b2  (
    .a({\picorv32_core/mem_rdata_latched [4],_al_u1627_o}),
    .b({_al_u1627_o,\picorv32_core/mem_rdata_latched [4]}),
    .c({_al_u1623_o,_al_u1623_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u1640_o,_al_u1640_o}),
    .mi({open_n28758,\picorv32_core/mem_rdata_latched [1]}),
    .q({open_n28765,\picorv32_core/decoded_rs2 [2]}));  // ../src/picorv32.v(1120)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*((~C*D)*~(0)*~(A)+(~C*D)*0*~(A)+~((~C*D))*0*A+(~C*D)*0*A))"),
    //.LUTF1("~B*~A*~C*D+B*~A*~C*D+~B*A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG0("(B*((~C*D)*~(1)*~(A)+(~C*D)*1*~(A)+~((~C*D))*1*A+(~C*D)*1*A))"),
    //.LUTG1("B*~A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*~A*~C*D+B*~A*~C*D+~B*A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000000),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b1000110010001000),
    .INIT_LUTG1(16'b1111111111111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg9_b3|_al_u1626  (
    .a({open_n28766,\picorv32_core/mem_rdata_latched$0$_placeOpt_3 }),
    .b({_al_u1627_o,\picorv32_core/mem_rdata_latched [1]}),
    .c({_al_u1623_o,_al_u1625_o}),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({_al_u1626_o,\picorv32_core/sel10_b3/B1_1 }),
    .e({_al_u1622_o,\picorv32_core/mem_rdata_latched [23]}),
    .f({open_n28782,_al_u1626_o}),
    .q({\picorv32_core/decoded_rs2 [3],open_n28786}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~((~A*~(C*B)))*~(D)+~0*(~A*~(C*B))*~(D)+~(~0)*(~A*~(C*B))*D+~0*(~A*~(C*B))*D)"),
    //.LUT1("~(~1*~((~A*~(C*B)))*~(D)+~1*(~A*~(C*B))*~(D)+~(~1)*(~A*~(C*B))*D+~1*(~A*~(C*B))*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110101000000000),
    .INIT_LUT1(16'b1110101011111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \picorv32_core/reg9_b4  (
    .a({_al_u1629_o,_al_u1629_o}),
    .b({_al_u1630_o,_al_u1630_o}),
    .c({\picorv32_core/n98_lutinv ,\picorv32_core/n98_lutinv }),
    .ce(\picorv32_core/n170 ),
    .clk(clk_pad),
    .d({\picorv32_core/n180 ,\picorv32_core/n180 }),
    .mi({open_n28797,\picorv32_core/mem_rdata_latched [24]}),
    .q({open_n28804,\picorv32_core/decoded_rs2 [4]}));  // ../src/picorv32.v(1120)
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u0|picorv32_core/sub0/ucin  (
    .a({\picorv32_core/pcpi_rs1$0$ ,1'b0}),
    .b({mem_la_wdata[0],open_n28805}),
    .f({\picorv32_core/n433 [0],open_n28825}),
    .fco(\picorv32_core/sub0/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u10|picorv32_core/sub0/u9  (
    .a({\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$9$ }),
    .b({\picorv32_core/pcpi_rs2$10$ ,\picorv32_core/pcpi_rs2$9$ }),
    .fci(\picorv32_core/sub0/c9 ),
    .f(\picorv32_core/n433 [10:9]),
    .fco(\picorv32_core/sub0/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u12|picorv32_core/sub0/u11  (
    .a({\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/pcpi_rs1$11$ }),
    .b({\picorv32_core/pcpi_rs2$12$ ,\picorv32_core/pcpi_rs2$11$ }),
    .fci(\picorv32_core/sub0/c11 ),
    .f(\picorv32_core/n433 [12:11]),
    .fco(\picorv32_core/sub0/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u14|picorv32_core/sub0/u13  (
    .a({\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$13$ }),
    .b({\picorv32_core/pcpi_rs2$14$ ,\picorv32_core/pcpi_rs2$13$ }),
    .fci(\picorv32_core/sub0/c13 ),
    .f(\picorv32_core/n433 [14:13]),
    .fco(\picorv32_core/sub0/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u16|picorv32_core/sub0/u15  (
    .a({\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/pcpi_rs1$15$ }),
    .b({\picorv32_core/pcpi_rs2$16$ ,\picorv32_core/pcpi_rs2$15$ }),
    .fci(\picorv32_core/sub0/c15 ),
    .f(\picorv32_core/n433 [16:15]),
    .fco(\picorv32_core/sub0/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u18|picorv32_core/sub0/u17  (
    .a({\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$17$ }),
    .b({\picorv32_core/pcpi_rs2$18$ ,\picorv32_core/pcpi_rs2$17$ }),
    .fci(\picorv32_core/sub0/c17 ),
    .f(\picorv32_core/n433 [18:17]),
    .fco(\picorv32_core/sub0/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u20|picorv32_core/sub0/u19  (
    .a({\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/pcpi_rs1$19$ }),
    .b({\picorv32_core/pcpi_rs2$20$ ,\picorv32_core/pcpi_rs2$19$ }),
    .fci(\picorv32_core/sub0/c19 ),
    .f(\picorv32_core/n433 [20:19]),
    .fco(\picorv32_core/sub0/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u22|picorv32_core/sub0/u21  (
    .a({\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs1$21$ }),
    .b({\picorv32_core/pcpi_rs2$22$ ,\picorv32_core/pcpi_rs2$21$ }),
    .fci(\picorv32_core/sub0/c21 ),
    .f(\picorv32_core/n433 [22:21]),
    .fco(\picorv32_core/sub0/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u24|picorv32_core/sub0/u23  (
    .a({\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/pcpi_rs1$23$ }),
    .b({\picorv32_core/pcpi_rs2$24$ ,\picorv32_core/pcpi_rs2$23$ }),
    .fci(\picorv32_core/sub0/c23 ),
    .f(\picorv32_core/n433 [24:23]),
    .fco(\picorv32_core/sub0/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u26|picorv32_core/sub0/u25  (
    .a({\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$25$ }),
    .b({\picorv32_core/pcpi_rs2$26$ ,\picorv32_core/pcpi_rs2$25$ }),
    .fci(\picorv32_core/sub0/c25 ),
    .f(\picorv32_core/n433 [26:25]),
    .fco(\picorv32_core/sub0/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u28|picorv32_core/sub0/u27  (
    .a({\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/pcpi_rs1$27$ }),
    .b({\picorv32_core/pcpi_rs2$28$ ,\picorv32_core/pcpi_rs2$27$ }),
    .fci(\picorv32_core/sub0/c27 ),
    .f(\picorv32_core/n433 [28:27]),
    .fco(\picorv32_core/sub0/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u2|picorv32_core/sub0/u1  (
    .a({\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$1$ }),
    .b(mem_la_wdata[2:1]),
    .fci(\picorv32_core/sub0/c1 ),
    .f(\picorv32_core/n433 [2:1]),
    .fco(\picorv32_core/sub0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u30|picorv32_core/sub0/u29  (
    .a({\picorv32_core/pcpi_rs1$30$ ,\picorv32_core/pcpi_rs1$29$ }),
    .b({\picorv32_core/pcpi_rs2$30$ ,\picorv32_core/pcpi_rs2$29$ }),
    .fci(\picorv32_core/sub0/c29 ),
    .f(\picorv32_core/n433 [30:29]),
    .fco(\picorv32_core/sub0/c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u31_al_u2577  (
    .a({open_n29094,\picorv32_core/pcpi_rs1$31$ }),
    .b({open_n29095,\picorv32_core/pcpi_rs2$31$ }),
    .fci(\picorv32_core/sub0/c31 ),
    .f({open_n29114,\picorv32_core/n433 [31]}));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u4|picorv32_core/sub0/u3  (
    .a({\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/pcpi_rs1$3$ }),
    .b(mem_la_wdata[4:3]),
    .fci(\picorv32_core/sub0/c3 ),
    .f(\picorv32_core/n433 [4:3]),
    .fco(\picorv32_core/sub0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u6|picorv32_core/sub0/u5  (
    .a({\picorv32_core/pcpi_rs1$6$ ,\picorv32_core/pcpi_rs1$5$ }),
    .b(mem_la_wdata[6:5]),
    .fci(\picorv32_core/sub0/c5 ),
    .f(\picorv32_core/n433 [6:5]),
    .fco(\picorv32_core/sub0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub0/u0|picorv32_core/sub0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub0/u8|picorv32_core/sub0/u7  (
    .a({\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/pcpi_rs1$7$ }),
    .b({\picorv32_core/pcpi_rs2$8$ ,mem_la_wdata[7]}),
    .fci(\picorv32_core/sub0/c7 ),
    .f(\picorv32_core/n433 [8:7]),
    .fco(\picorv32_core/sub0/c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub1/u0|picorv32_core/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub1/u0|picorv32_core/sub1/ucin  (
    .a({\picorv32_core/reg_sh [0],1'b0}),
    .b({1'b0,open_n29186}),
    .f({\picorv32_core/n559 [0],open_n29206}),
    .fco(\picorv32_core/sub1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub1/u0|picorv32_core/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub1/u2|picorv32_core/sub1/u1  (
    .a(\picorv32_core/reg_sh [2:1]),
    .b(2'b10),
    .fci(\picorv32_core/sub1/c1 ),
    .f(\picorv32_core/n559 [2:1]),
    .fco(\picorv32_core/sub1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub1/u0|picorv32_core/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub1/u4|picorv32_core/sub1/u3  (
    .a(\picorv32_core/reg_sh [4:3]),
    .b(2'b00),
    .fci(\picorv32_core/sub1/c3 ),
    .f(\picorv32_core/n559 [4:3]));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub2/u0|picorv32_core/sub2/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub2/u0|picorv32_core/sub2/ucin  (
    .a({\picorv32_core/reg_sh [0],1'b0}),
    .b({1'b1,open_n29256}),
    .f({\picorv32_core/n564 [0],open_n29276}),
    .fco(\picorv32_core/sub2/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub2/u0|picorv32_core/sub2/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub2/u2|picorv32_core/sub2/u1  (
    .a(\picorv32_core/reg_sh [2:1]),
    .b(2'b00),
    .fci(\picorv32_core/sub2/c1 ),
    .f(\picorv32_core/n564 [2:1]),
    .fco(\picorv32_core/sub2/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("picorv32_core/sub2/u0|picorv32_core/sub2/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \picorv32_core/sub2/u4|picorv32_core/sub2/u3  (
    .a(\picorv32_core/reg_sh [4:3]),
    .b(2'b00),
    .fci(\picorv32_core/sub2/c3 ),
    .f(\picorv32_core/n564 [4:3]));
  // ../src/top.v(42)
  // ../src/top.v(42)
  EG_PHY_LSLICE #(
    //.LUTF0("(A@D)"),
    //.LUTF1("(~A)"),
    //.LUTG0("(A@D)"),
    //.LUTG1("(~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010110101010),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0101010110101010),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \reg0_b0|reg0_b1  (
    .a({initial_reset[0],initial_reset[1]}),
    .ce(\eq0/or_xor_i0$0$_i1$0$_o_o ),
    .clk(clk_pad),
    .d({open_n29330,initial_reset[0]}),
    .q({initial_reset[0],initial_reset[1]}));  // ../src/top.v(42)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P10"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("SET"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTRSTMUX("INV"),
    .OUTSCLKMUX("CLK"),
    .SRMODE("ASYNC"),
    .TSMUX("0"))
    reg1_b0_DO (
    .ce(n16),
    .do({open_n29353,open_n29354,open_n29355,n17[0]}),
    .osclk(clk_pad),
    .rst(resetn_placeOpt_4),
    .opad(out_byte[0]));  // ../src/top.v(128)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("SET"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTRSTMUX("INV"),
    .OUTSCLKMUX("CLK"),
    .SRMODE("ASYNC"),
    .TSMUX("0"))
    reg1_b1_DO (
    .ce(n16),
    .do({open_n29367,open_n29368,open_n29369,n17[1]}),
    .osclk(clk_pad),
    .rst(resetn_placeOpt_6),
    .opad(out_byte[1]));  // ../src/top.v(128)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("SET"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTRSTMUX("INV"),
    .OUTSCLKMUX("CLK"),
    .SRMODE("ASYNC"),
    .TSMUX("0"))
    reg1_b2_DO (
    .ce(n16),
    .do({open_n29381,open_n29382,open_n29383,n17[2]}),
    .osclk(clk_pad),
    .rst(resetn_placeOpt_6),
    .opad(out_byte[2]));  // ../src/top.v(128)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("SET"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTRSTMUX("INV"),
    .OUTSCLKMUX("CLK"),
    .SRMODE("ASYNC"),
    .TSMUX("0"))
    reg1_b3_DO (
    .ce(n16),
    .do({open_n29395,open_n29396,open_n29397,n17[3]}),
    .osclk(clk_pad),
    .rst(resetn_placeOpt_6),
    .opad(out_byte[3]));  // ../src/top.v(128)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("SET"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTRSTMUX("INV"),
    .OUTSCLKMUX("CLK"),
    .SRMODE("ASYNC"),
    .TSMUX("0"))
    reg1_b4_DO (
    .ce(n16),
    .do({open_n29409,open_n29410,open_n29411,n17[4]}),
    .osclk(clk_pad),
    .rst(resetn_placeOpt_6),
    .opad(out_byte[4]));  // ../src/top.v(128)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P17"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("SET"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTRSTMUX("INV"),
    .OUTSCLKMUX("CLK"),
    .SRMODE("ASYNC"),
    .TSMUX("0"))
    reg1_b5_DO (
    .ce(n16),
    .do({open_n29423,open_n29424,open_n29425,n17[5]}),
    .osclk(clk_pad),
    .rst(resetn_placeOpt_1),
    .opad(out_byte[5]));  // ../src/top.v(128)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P19"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("SET"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTRSTMUX("INV"),
    .OUTSCLKMUX("CLK"),
    .SRMODE("ASYNC"),
    .TSMUX("0"))
    reg1_b6_DO (
    .ce(n16),
    .do({open_n29437,open_n29438,open_n29439,n17[6]}),
    .osclk(clk_pad),
    .rst(resetn_placeOpt_3),
    .opad(out_byte[6]));  // ../src/top.v(128)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P23"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("SET"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTRSTMUX("INV"),
    .OUTSCLKMUX("CLK"),
    .SRMODE("ASYNC"),
    .TSMUX("0"))
    reg1_b7_DO (
    .ce(n16),
    .do({open_n29451,open_n29452,open_n29453,n17[7]}),
    .osclk(clk_pad),
    .rst(resetn_placeOpt_11),
    .opad(out_byte[7]));  // ../src/top.v(128)
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u0|uart/add0/ucin  (
    .a({\uart/uart_counter [0],1'b0}),
    .b({1'b1,open_n29465}),
    .f({\uart/n5 [0],open_n29485}),
    .fco(\uart/add0/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u10|uart/add0/u9  (
    .a(\uart/uart_counter [10:9]),
    .b(2'b00),
    .fci(\uart/add0/c9 ),
    .f(\uart/n5 [10:9]),
    .fco(\uart/add0/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u12|uart/add0/u11  (
    .a({1'b0,\uart/uart_counter [11]}),
    .b({\uart/uart_counter [12],1'b0}),
    .fci(\uart/add0/c11 ),
    .f(\uart/n5 [12:11]),
    .fco(\uart/add0/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u14|uart/add0/u13  (
    .a(2'b00),
    .b(\uart/uart_counter [14:13]),
    .fci(\uart/add0/c13 ),
    .f(\uart/n5 [14:13]),
    .fco(\uart/add0/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u16|uart/add0/u15  (
    .a({\uart/uart_counter [16],1'b0}),
    .b({1'b0,\uart/uart_counter [15]}),
    .fci(\uart/add0/c15 ),
    .f(\uart/n5 [16:15]),
    .fco(\uart/add0/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u18|uart/add0/u17  (
    .a({1'b0,\uart/uart_counter [17]}),
    .b({\uart/uart_counter [18],1'b0}),
    .fci(\uart/add0/c17 ),
    .f(\uart/n5 [18:17]),
    .fco(\uart/add0/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u20|uart/add0/u19  (
    .a(\uart/uart_counter [20:19]),
    .b(2'b00),
    .fci(\uart/add0/c19 ),
    .f(\uart/n5 [20:19]),
    .fco(\uart/add0/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u22|uart/add0/u21  (
    .a({\uart/uart_counter [22],1'b0}),
    .b({1'b0,\uart/uart_counter [21]}),
    .fci(\uart/add0/c21 ),
    .f(\uart/n5 [22:21]),
    .fco(\uart/add0/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u24|uart/add0/u23  (
    .a(\uart/uart_counter [24:23]),
    .b(2'b00),
    .fci(\uart/add0/c23 ),
    .f(\uart/n5 [24:23]),
    .fco(\uart/add0/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u26|uart/add0/u25  (
    .a({\uart/uart_counter [26],1'b0}),
    .b({1'b0,\uart/uart_counter [25]}),
    .fci(\uart/add0/c25 ),
    .f(\uart/n5 [26:25]),
    .fco(\uart/add0/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u28|uart/add0/u27  (
    .a({\uart/uart_counter [28],1'b0}),
    .b({1'b0,\uart/uart_counter [27]}),
    .fci(\uart/add0/c27 ),
    .f(\uart/n5 [28:27]),
    .fco(\uart/add0/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u2|uart/add0/u1  (
    .a({\uart/uart_counter [2],1'b0}),
    .b({1'b0,\uart/uart_counter [1]}),
    .fci(\uart/add0/c1 ),
    .f(\uart/n5 [2:1]),
    .fco(\uart/add0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u30|uart/add0/u29  (
    .a(2'b00),
    .b(\uart/uart_counter [30:29]),
    .fci(\uart/add0/c29 ),
    .f(\uart/n5 [30:29]),
    .fco(\uart/add0/c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u31_al_u2578  (
    .a({open_n29754,\uart/uart_counter [31]}),
    .b({open_n29755,1'b0}),
    .fci(\uart/add0/c31 ),
    .f({open_n29774,\uart/n5 [31]}));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u4|uart/add0/u3  (
    .a(2'b00),
    .b(\uart/uart_counter [4:3]),
    .fci(\uart/add0/c3 ),
    .f(\uart/n5 [4:3]),
    .fco(\uart/add0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u6|uart/add0/u5  (
    .a({1'b0,\uart/uart_counter [5]}),
    .b({\uart/uart_counter [6],1'b0}),
    .fci(\uart/add0/c5 ),
    .f(\uart/n5 [6:5]),
    .fco(\uart/add0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add0/u0|uart/add0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add0/u8|uart/add0/u7  (
    .a(2'b00),
    .b(\uart/uart_counter [8:7]),
    .fci(\uart/add0/c7 ),
    .f(\uart/n5 [8:7]),
    .fco(\uart/add0/c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add1/u0|uart/add1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add1/u0|uart/add1/ucin  (
    .a({\uart/uart_status_txd [0],1'b0}),
    .b({1'b1,open_n29846}),
    .f({\uart/n35 [0],open_n29866}),
    .fco(\uart/add1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add1/u0|uart/add1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add1/u2|uart/add1/u1  (
    .a({1'b0,\uart/uart_status_txd [1]}),
    .b({\uart/uart_status_txd [2],1'b0}),
    .fci(\uart/add1/c1 ),
    .f(\uart/n35 [2:1]),
    .fco(\uart/add1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add1/u0|uart/add1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add1/u3_al_u2579  (
    .a({open_n29893,1'b0}),
    .b({open_n29894,\uart/uart_status_txd [3]}),
    .fci(\uart/add1/c3 ),
    .f({open_n29913,\uart/n35 [3]}));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add2/u0|uart/add2/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add2/u0|uart/add2/ucin  (
    .a({\uart/uart_smp_rx [0],1'b0}),
    .b({1'b1,open_n29919}),
    .f({\uart/n49 [0],open_n29939}),
    .fco(\uart/add2/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add2/u0|uart/add2/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add2/u2|uart/add2/u1  (
    .a(\uart/uart_smp_rx [2:1]),
    .b(2'b00),
    .fci(\uart/add2/c1 ),
    .f(\uart/n49 [2:1]),
    .fco(\uart/add2/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add2/u0|uart/add2/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add2/u3_al_u2580  (
    .a({open_n29966,1'b0}),
    .b({open_n29967,\uart/uart_smp_rx [3]}),
    .fci(\uart/add2/c3 ),
    .f({open_n29986,\uart/n49 [3]}));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add3/u0|uart/add3/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add3/u0|uart/add3/ucin  (
    .a({\uart/uart_status_rxd [0],1'b0}),
    .b({1'b1,open_n29992}),
    .f({\uart/n77 [0],open_n30012}),
    .fco(\uart/add3/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add3/u0|uart/add3/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add3/u2|uart/add3/u1  (
    .a({1'b0,\uart/uart_status_rxd [1]}),
    .b({\uart/uart_status_rxd [2],1'b0}),
    .fci(\uart/add3/c1 ),
    .f(\uart/n77 [2:1]),
    .fco(\uart/add3/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/add3/u0|uart/add3/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \uart/add3/u3_al_u2581  (
    .a({open_n30039,1'b0}),
    .b({open_n30040,\uart/uart_status_rxd [3]}),
    .fci(\uart/add3/c3 ),
    .f({open_n30059,\uart/n77 [3]}));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_0|uart/lt0_cin  (
    .a({\uart/uart_bsrr [0],1'b1}),
    .b({\uart/uart_counter [0],open_n30065}),
    .fco(\uart/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_10|uart/lt0_9  (
    .a(\uart/uart_bsrr [10:9]),
    .b(\uart/uart_counter [10:9]),
    .fci(\uart/lt0_c9 ),
    .fco(\uart/lt0_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_12|uart/lt0_11  (
    .a(\uart/uart_bsrr [12:11]),
    .b(\uart/uart_counter [12:11]),
    .fci(\uart/lt0_c11 ),
    .fco(\uart/lt0_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_14|uart/lt0_13  (
    .a(\uart/uart_bsrr [14:13]),
    .b(\uart/uart_counter [14:13]),
    .fci(\uart/lt0_c13 ),
    .fco(\uart/lt0_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_16|uart/lt0_15  (
    .a(\uart/uart_bsrr [16:15]),
    .b(\uart/uart_counter [16:15]),
    .fci(\uart/lt0_c15 ),
    .fco(\uart/lt0_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_18|uart/lt0_17  (
    .a(\uart/uart_bsrr [18:17]),
    .b(\uart/uart_counter [18:17]),
    .fci(\uart/lt0_c17 ),
    .fco(\uart/lt0_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_20|uart/lt0_19  (
    .a(\uart/uart_bsrr [20:19]),
    .b(\uart/uart_counter [20:19]),
    .fci(\uart/lt0_c19 ),
    .fco(\uart/lt0_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_22|uart/lt0_21  (
    .a(\uart/uart_bsrr [22:21]),
    .b(\uart/uart_counter [22:21]),
    .fci(\uart/lt0_c21 ),
    .fco(\uart/lt0_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_24|uart/lt0_23  (
    .a(\uart/uart_bsrr [24:23]),
    .b(\uart/uart_counter [24:23]),
    .fci(\uart/lt0_c23 ),
    .fco(\uart/lt0_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_26|uart/lt0_25  (
    .a(\uart/uart_bsrr [26:25]),
    .b(\uart/uart_counter [26:25]),
    .fci(\uart/lt0_c25 ),
    .fco(\uart/lt0_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_28|uart/lt0_27  (
    .a(\uart/uart_bsrr [28:27]),
    .b(\uart/uart_counter [28:27]),
    .fci(\uart/lt0_c27 ),
    .fco(\uart/lt0_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_2|uart/lt0_1  (
    .a(\uart/uart_bsrr [2:1]),
    .b(\uart/uart_counter [2:1]),
    .fci(\uart/lt0_c1 ),
    .fco(\uart/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_30|uart/lt0_29  (
    .a(\uart/uart_bsrr [30:29]),
    .b(\uart/uart_counter [30:29]),
    .fci(\uart/lt0_c29 ),
    .fco(\uart/lt0_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_4|uart/lt0_3  (
    .a(\uart/uart_bsrr [4:3]),
    .b(\uart/uart_counter [4:3]),
    .fci(\uart/lt0_c3 ),
    .fco(\uart/lt0_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_6|uart/lt0_5  (
    .a(\uart/uart_bsrr [6:5]),
    .b(\uart/uart_counter [6:5]),
    .fci(\uart/lt0_c5 ),
    .fco(\uart/lt0_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \uart/lt0_8|uart/lt0_7  (
    .a(\uart/uart_bsrr [8:7]),
    .b(\uart/uart_counter [8:7]),
    .fci(\uart/lt0_c7 ),
    .fco(\uart/lt0_c9 ));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(0*~A)*~(~B*C))"),
    //.LUT1("~(~D*~(1*~A)*~(~B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1111111101110101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg0_b0  (
    .a({_al_u812_o,_al_u812_o}),
    .b({_al_u894_o,_al_u894_o}),
    .c({_al_u892_o,_al_u892_o}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({_al_u893_o,_al_u893_o}),
    .mi({open_n30461,\uart/uart_bsrr [0]}),
    .sr(resetn),
    .q({open_n30467,uart_do[0]}));  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(0*~A)*~(~B*C))"),
    //.LUT1("~(~D*~(1*~A)*~(~B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1111111101110101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg0_b1  (
    .a({_al_u812_o,_al_u812_o}),
    .b({_al_u817_o,_al_u817_o}),
    .c({_al_u815_o,_al_u815_o}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({_al_u816_o,_al_u816_o}),
    .mi({open_n30478,\uart/uart_bsrr [1]}),
    .sr(resetn),
    .q({open_n30484,uart_do[1]}));  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(0*~A)*~(~B*C))"),
    //.LUT1("~(~D*~(1*~A)*~(~B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1111111101110101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg0_b2  (
    .a({_al_u812_o,_al_u812_o}),
    .b({_al_u813_o,_al_u813_o}),
    .c({_al_u810_o,_al_u810_o}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({_al_u811_o,_al_u811_o}),
    .mi({open_n30495,\uart/uart_bsrr [2]}),
    .sr(resetn),
    .q({open_n30501,uart_do[2]}));  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*C*~(A)*~(0)+~(D)*~(B)*~(C)*A*~(0)+~(D)*~(B)*C*A*~(0)+D*~(B)*C*A*~(0)+~(D)*B*~(C)*~(A)*0+D*~(B)*C*~(A)*0+~(D)*B*C*~(A)*0+~(D)*~(B)*~(C)*A*0+~(D)*B*~(C)*A*0+~(D)*~(B)*C*A*0+D*~(B)*C*A*0+~(D)*B*C*A*0)"),
    //.LUT1("(C*~(B)*A*~(D)*~(1)+~(C)*~(B)*~(A)*D*~(1)+~(C)*~(B)*A*D*~(1)+C*~(B)*A*D*~(1)+~(C)*B*~(A)*~(D)*1+C*~(B)*A*~(D)*1+~(C)*B*A*~(D)*1+~(C)*~(B)*~(A)*D*1+~(C)*B*~(A)*D*1+~(C)*~(B)*A*D*1+C*~(B)*A*D*1+~(C)*B*A*D*1)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000000100010),
    .INIT_LUT1(16'b0010111100101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg0_b5  (
    .a({\uart/uart_bsrr [5],\uart/uart_odr [5]}),
    .b({mem_la_addr[2],mem_la_addr[2]}),
    .c({mem_la_addr[3],\uart/uart_bsrr [5]}),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({\uart/uart_odr [5],mem_la_addr[3]}),
    .mi({open_n30512,\uart/uart_idr [5]}),
    .sr(resetn),
    .q({open_n30518,uart_do[5]}));  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C)*B*~(A)*~(0)+~(D)*~(C)*~(B)*A*~(0)+~(D)*~(C)*B*A*~(0)+D*~(C)*B*A*~(0)+~(D)*C*~(B)*~(A)*0+D*~(C)*B*~(A)*0+~(D)*C*B*~(A)*0+~(D)*~(C)*~(B)*A*0+~(D)*C*~(B)*A*0+~(D)*~(C)*B*A*0+D*~(C)*B*A*0+~(D)*C*B*A*0)"),
    //.LUT1("(C*~(D)*A*~(B)*~(1)+~(C)*~(D)*~(A)*B*~(1)+~(C)*~(D)*A*B*~(1)+C*~(D)*A*B*~(1)+~(C)*D*~(A)*~(B)*1+C*~(D)*A*~(B)*1+~(C)*D*A*~(B)*1+~(C)*~(D)*~(A)*B*1+~(C)*D*~(A)*B*1+~(C)*~(D)*A*B*1+C*~(D)*A*B*1+~(C)*D*A*B*1)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b0000111110101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg0_b6  (
    .a({\uart/uart_bsrr [6],\uart/uart_odr [6]}),
    .b({\uart/uart_odr [6],\uart/uart_bsrr [6]}),
    .c(mem_la_addr[3:2]),
    .ce(\uart/mux14_b0_sel_is_1_o ),
    .clk(clk_pad),
    .d({mem_la_addr[2],mem_la_addr[3]}),
    .mi({open_n30529,\uart/uart_idr [6]}),
    .sr(resetn),
    .q({open_n30535,uart_do[6]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000001010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg10_b0|uart/reg10_b1  (
    .a({\uart/n4 [1],open_n30536}),
    .c({open_n30539,\uart/uart_op_clock }),
    .ce(\uart/n2 ),
    .clk(clk_pad),
    .d({\uart/uart_op_clock_by_3_c [1],\uart/n4 [1]}),
    .mi({open_n30550,\uart/n4 [1]}),
    .sr(resetn_placeOpt_5),
    .f({open_n30551,_al_u1076_o}),
    .q({\uart/n4 [1],\uart/uart_op_clock_by_3_c [1]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~D)"),
    //.LUTF1("(B*~D)"),
    //.LUTG0("(B*~D)"),
    //.LUTG1("(B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001100),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b0000000011001100),
    .INIT_LUTG1(16'b0000000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b0|uart/reg1_b9  (
    .b({\uart/n5 [0],\uart/n5 [9]}),
    .clk(clk_pad),
    .d({\uart/n2 ,\uart/n2 }),
    .sr(resetn_placeOpt_2),
    .q({\uart/uart_counter [0],\uart/uart_counter [9]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~C)"),
    //.LUT1("(D*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110000001100),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b10|uart/reg1_b8  (
    .b({\uart/n2 ,\uart/n5 [8]}),
    .c({open_n30583,\uart/n2 }),
    .clk(clk_pad),
    .d({\uart/n5 [10],open_n30585}),
    .sr(resetn_placeOpt_2),
    .q({\uart/uart_counter [10],\uart/uart_counter [8]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A)"),
    //.LUT1("(C*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000001010000),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b11|uart/reg1_b7  (
    .a({\uart/n2 ,\uart/n2 }),
    .c({\uart/n5 [11],\uart/n5 [7]}),
    .clk(clk_pad),
    .sr(resetn_placeOpt_2),
    .q({\uart/uart_counter [11],\uart/uart_counter [7]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("0"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*~C*B*D+A*~C*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b12|uart/reg1_b6  (
    .c({\uart/n2 ,\uart/n5 [6]}),
    .clk(clk_pad),
    .d({open_n30630,\uart/n2 }),
    .e({\uart/n5 [12],open_n30631}),
    .sr(resetn_placeOpt_2),
    .q({\uart/uart_counter [12],\uart/uart_counter [6]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A)"),
    //.LUTF1("(D*~C)"),
    //.LUTG0("(C*~A)"),
    //.LUTG1("(D*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0101000001010000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b13|uart/reg1_b5  (
    .a({open_n30651,\uart/n2 }),
    .c({\uart/n2 ,\uart/n5 [5]}),
    .clk(clk_pad),
    .d({\uart/n5 [13],open_n30655}),
    .sr(resetn_placeOpt_2),
    .q({\uart/uart_counter [13],\uart/uart_counter [5]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A)"),
    //.LUT1("(C*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000001010000),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b14|uart/reg1_b4  (
    .a({\uart/n2 ,\uart/n2 }),
    .c({\uart/n5 [14],\uart/n5 [4]}),
    .clk(clk_pad),
    .sr(resetn_placeOpt_2),
    .q({\uart/uart_counter [14],\uart/uart_counter [4]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A)"),
    //.LUT1("(C*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000001010000),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b15|uart/reg1_b31  (
    .a({\uart/n2 ,\uart/n2 }),
    .c({\uart/n5 [15],\uart/n5 [31]}),
    .clk(clk_pad),
    .sr(resetn_placeOpt_5),
    .q({\uart/uart_counter [15],\uart/uart_counter [31]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(A*~C)"),
    //.LUTG0("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C"),
    //.LUTG1("(A*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000101000001010),
    .INIT_LUTG0(16'b0000111100001111),
    .INIT_LUTG1(16'b0000101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b16|uart/reg1_b30  (
    .a({\uart/n5 [16],open_n30721}),
    .c({\uart/n2 ,\uart/n2 }),
    .clk(clk_pad),
    .e({open_n30727,\uart/n5 [30]}),
    .sr(resetn_placeOpt_5),
    .q({\uart/uart_counter [16],\uart/uart_counter [30]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b17|uart/reg1_b3  (
    .b({\uart/n5 [17],open_n30749}),
    .c({open_n30750,\uart/n5 [3]}),
    .clk(clk_pad),
    .d({\uart/n2 ,\uart/n2 }),
    .sr(resetn_placeOpt_2),
    .q({\uart/uart_counter [17],\uart/uart_counter [3]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A)"),
    //.LUT1("(C*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000001010000),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b18|uart/reg1_b29  (
    .a({\uart/n2 ,\uart/n2 }),
    .c({\uart/n5 [18],\uart/n5 [29]}),
    .clk(clk_pad),
    .sr(resetn_placeOpt_5),
    .q({\uart/uart_counter [18],\uart/uart_counter [29]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~B)"),
    //.LUT1("(D*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001000100010),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b19|uart/reg1_b28  (
    .a({open_n30795,\uart/n5 [28]}),
    .b({\uart/n2 ,\uart/n2 }),
    .clk(clk_pad),
    .d({\uart/n5 [19],open_n30799}),
    .sr(resetn_placeOpt_5),
    .q({\uart/uart_counter [19],\uart/uart_counter [28]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A)"),
    //.LUTF1("(D*~C)"),
    //.LUTG0("(C*~A)"),
    //.LUTG1("(D*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0101000001010000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b1|uart/reg1_b27  (
    .a({open_n30817,\uart/n2 }),
    .c({\uart/n2 ,\uart/n5 [27]}),
    .clk(clk_pad),
    .d({\uart/n5 [1],open_n30821}),
    .sr(resetn_placeOpt_2),
    .q({\uart/uart_counter [1],\uart/uart_counter [27]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(B*~D)"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG1("(B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b0000000011111111),
    .INIT_LUTG1(16'b0000000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b20|uart/reg1_b26  (
    .b({\uart/n5 [20],open_n30845}),
    .clk(clk_pad),
    .d({\uart/n2 ,\uart/n2 }),
    .e({open_n30849,\uart/n5 [26]}),
    .sr(resetn_placeOpt_5),
    .q({\uart/uart_counter [20],\uart/uart_counter [26]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~C)"),
    //.LUT1("(B*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110000001100),
    .INIT_LUT1(16'b0000110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b21|uart/reg1_b25  (
    .b({\uart/n5 [21],\uart/n5 [25]}),
    .c({\uart/n2 ,\uart/n2 }),
    .clk(clk_pad),
    .sr(resetn_placeOpt_5),
    .q({\uart/uart_counter [21],\uart/uart_counter [25]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B)"),
    //.LUT1("(D*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000000110000),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b22|uart/reg1_b24  (
    .b({\uart/n2 ,\uart/n2 }),
    .c({open_n30893,\uart/n5 [24]}),
    .clk(clk_pad),
    .d({\uart/n5 [22],open_n30895}),
    .sr(resetn_placeOpt_5),
    .q({\uart/uart_counter [22],\uart/uart_counter [24]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~D)"),
    //.LUTF1("0"),
    //.LUTG0("(B*~D)"),
    //.LUTG1("~D*~B*~C*~A+~D*B*~C*~A+~D*~B*C*~A+~D*B*C*~A+~D*~B*~C*A+~D*B*~C*A+~D*~B*C*A+~D*B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001100),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000011001100),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg1_b2|uart/reg1_b23  (
    .b({open_n30915,\uart/n5 [23]}),
    .clk(clk_pad),
    .d({\uart/n2 ,\uart/n2 }),
    .e({\uart/n5 [2],open_n30919}),
    .sr(resetn_placeOpt_2),
    .q({\uart/uart_counter [2],\uart/uart_counter [23]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("~B*~D*~C*A+B*~D*~C*A+~B*~D*C*A+B*~D*C*A"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("~B*D*~C*~A+B*D*~C*~A+~B*D*C*~A+B*D*C*~A+~B*~D*~C*A+B*~D*~C*A+~B*D*~C*A+B*D*~C*A+~B*~D*C*A+B*~D*C*A+~B*D*C*A+B*D*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b0000000010101010),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b1111111110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg2_b11|uart/reg2_b3  (
    .a({\picorv32_core/pcpi_rs2$11$ ,_al_u826_o}),
    .b({open_n30939,_al_u827_o}),
    .c({open_n30940,_al_u828_o}),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_wordsize [1],\picorv32_core/pcpi_rs1$3$ }),
    .e({mem_la_wdata[3],mem_la_wdata[3]}),
    .mi({open_n30942,mem_la_wdata[3]}),
    .sr(resetn_placeOpt_2),
    .f({mem_la_wdata[11],_al_u873_o}),
    .q({\uart/uart_bsrr [11],\uart/uart_bsrr [3]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B)*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A"),
    //.LUTG0("(A*~(B)*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000100100000),
    .INIT_LUTF1(16'b0000101000001010),
    .INIT_LUTG0(16'b0111010101100100),
    .INIT_LUTG1(16'b1111101011111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg2_b12|uart/reg2_b28  (
    .a({\picorv32_core/pcpi_rs2$12$ ,\picorv32_core/mem_wordsize [0]}),
    .b({open_n30957,\picorv32_core/mem_wordsize [1]}),
    .c({\picorv32_core/mem_wordsize [1],\picorv32_core/pcpi_rs2$12$ }),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({open_n30958,\picorv32_core/pcpi_rs2$28$ }),
    .e({mem_la_wdata[4],mem_la_wdata[4]}),
    .sr(resetn_placeOpt_12),
    .f({mem_la_wdata[12],mem_la_wdata[28]}),
    .q({\uart/uart_bsrr [12],\uart/uart_bsrr [28]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("A*~D*~C*B+A*D*~C*B+A*~D*C*B+A*D*C*B"),
    //.LUTG0("(~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+A*~D*~C*B+A*D*~C*B+A*~D*C*B+A*D*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100000000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b0011111101110111),
    .INIT_LUTG1(16'b1011101110111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg2_b13|uart/reg2_b5  (
    .a({mem_la_wdata[5],_al_u826_o}),
    .b({\picorv32_core/mem_wordsize [1],_al_u827_o}),
    .c({open_n30976,_al_u828_o}),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({open_n30977,\picorv32_core/pcpi_rs1$5$ }),
    .e({\picorv32_core/pcpi_rs2$13$ ,mem_la_wdata[5]}),
    .mi({open_n30979,mem_la_wdata[5]}),
    .sr(resetn_placeOpt_2),
    .f({mem_la_wdata[13],_al_u881_o}),
    .q({\uart/uart_bsrr [13],\uart/uart_bsrr [5]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B)*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(A*~(B)*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000100100000),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b0111010101100100),
    .INIT_LUTG1(16'b1111111111001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg2_b14|uart/reg2_b30  (
    .a({open_n30994,\picorv32_core/mem_wordsize [0]}),
    .b({\picorv32_core/pcpi_rs2$14$ ,\picorv32_core/mem_wordsize [1]}),
    .c({open_n30995,\picorv32_core/pcpi_rs2$14$ }),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_wordsize [1],\picorv32_core/pcpi_rs2$30$ }),
    .e({mem_la_wdata[6],mem_la_wdata[6]}),
    .sr(resetn_placeOpt_12),
    .f({mem_la_wdata[14],mem_la_wdata[30]}),
    .q({\uart/uart_bsrr [14],\uart/uart_bsrr [30]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B)*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("C*~B*~A*~D+C*B*~A*~D+C*~B*A*~D+C*B*A*~D"),
    //.LUTG0("(A*~(B)*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("C*~B*~A*~D+C*B*~A*~D+C*~B*A*~D+C*B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000100100000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0111010101100100),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg2_b15|uart/reg2_b31  (
    .a({open_n31013,\picorv32_core/mem_wordsize [0]}),
    .b({open_n31014,\picorv32_core/mem_wordsize [1]}),
    .c({\picorv32_core/pcpi_rs2$15$ ,\picorv32_core/pcpi_rs2$15$ }),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\picorv32_core/mem_wordsize [1],\picorv32_core/pcpi_rs2$31$ }),
    .e({mem_la_wdata[7],mem_la_wdata[7]}),
    .sr(resetn_placeOpt_12),
    .f({mem_la_wdata[15],mem_la_wdata[31]}),
    .q({\uart/uart_bsrr [15],\uart/uart_bsrr [31]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100101011001010),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg2_b16|uart/reg2_b22  (
    .a({open_n31032,mem_la_wdata[6]}),
    .b({\picorv32_core/n734_lutinv ,\picorv32_core/pcpi_rs2$22$ }),
    .c({mem_la_wdata[0],\picorv32_core/n734_lutinv }),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\picorv32_core/pcpi_rs2$16$ ,open_n31033}),
    .sr(resetn_placeOpt_13),
    .f({mem_la_wdata[16],mem_la_wdata[22]}),
    .q({\uart/uart_bsrr [16],\uart/uart_bsrr [22]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*A*~D*C+B*A*~D*C+~B*A*D*C+B*A*D*C"),
    //.LUTF1("~D*~C*B*A+D*~C*B*A+~D*C*B*A+D*C*B*A"),
    //.LUTG0("~B*~A*~D*~C+B*~A*~D*~C+~B*A*~D*~C+B*A*~D*~C+~B*~A*D*~C+B*~A*D*~C+~B*A*D*~C+B*A*D*~C+~B*A*~D*C+B*A*~D*C+~B*A*D*C+B*A*D*C"),
    //.LUTG1("~D*~C*~B*~A+D*~C*~B*~A+~D*C*~B*~A+D*C*~B*~A+~D*~C*~B*A+D*~C*~B*A+~D*C*~B*A+D*C*~B*A+~D*~C*B*A+D*~C*B*A+~D*C*B*A+D*C*B*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010000010100000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1010111110101111),
    .INIT_LUTG1(16'b1011101110111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg2_b17|uart/reg2_b9  (
    .a({\picorv32_core/pcpi_rs2$17$ ,mem_la_wdata[1]}),
    .b({\picorv32_core/n734_lutinv ,open_n31049}),
    .c({open_n31050,\picorv32_core/mem_wordsize [1]}),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .e({mem_la_wdata[1],\picorv32_core/pcpi_rs2$9$ }),
    .sr(resetn),
    .f({mem_la_wdata[17],mem_la_wdata[9]}),
    .q({\uart/uart_bsrr [17],\uart/uart_bsrr [9]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110001011100010),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg2_b18|uart/reg2_b10  (
    .a({open_n31070,\picorv32_core/pcpi_rs2$10$ }),
    .b({\picorv32_core/n734_lutinv ,\picorv32_core/mem_wordsize [1]}),
    .c({mem_la_wdata[2],mem_la_wdata[2]}),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\picorv32_core/pcpi_rs2$18$ ,open_n31071}),
    .sr(resetn_placeOpt_12),
    .f({mem_la_wdata[18],mem_la_wdata[10]}),
    .q({\uart/uart_bsrr [18],\uart/uart_bsrr [10]}));  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*~(B)*~(C)*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUT1("(~(C)*B*A*~(D)*~(1)+~(C)*~(B)*~(A)*D*~(1)+~(C)*~(B)*A*D*~(1)+~(C)*B*A*D*~(1)+C*~(B)*~(A)*~(D)*1+C*~(B)*A*~(D)*1+~(C)*B*A*~(D)*1+~(C)*~(B)*~(A)*D*1+C*~(B)*~(A)*D*1+~(C)*~(B)*A*D*1+C*~(B)*A*D*1+~(C)*B*A*D*1)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0011101100111000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg2_b25  (
    .a({mem_la_wdata[1],\picorv32_core/mem_wordsize [0]}),
    .b({\picorv32_core/mem_wordsize [1],\picorv32_core/mem_wordsize [1]}),
    .c({\picorv32_core/mem_wordsize [0],mem_la_wdata[1]}),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\picorv32_core/pcpi_rs2$25$ ,\picorv32_core/pcpi_rs2$25$ }),
    .mi({open_n31097,\picorv32_core/pcpi_rs2$9$ }),
    .sr(resetn_placeOpt_13),
    .fx({open_n31101,mem_la_wdata[25]}),
    .q({open_n31102,\uart/uart_bsrr [25]}));  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*C*~(D)*~(0)+~(A)*B*~(C)*D*~(0)+A*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUT1("(C*~(B)*A*~(D)*~(1)+~(C)*B*~(A)*D*~(1)+C*~(B)*A*D*~(1)+~(C)*B*A*D*~(1)+~(C)*~(B)*~(A)*~(D)*1+~(C)*~(B)*A*~(D)*1+C*~(B)*A*~(D)*1+~(C)*~(B)*~(A)*D*1+~(C)*B*~(A)*D*1+~(C)*~(B)*A*D*1+C*~(B)*A*D*1+~(C)*B*A*D*1)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0110010000100000),
    .INIT_LUT1(16'b0010111100100011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg2_b26  (
    .a({\picorv32_core/pcpi_rs2$10$ ,\picorv32_core/mem_wordsize [0]}),
    .b({\picorv32_core/mem_wordsize [1],\picorv32_core/mem_wordsize [1]}),
    .c({\picorv32_core/mem_wordsize [0],\picorv32_core/pcpi_rs2$10$ }),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({mem_la_wdata[2],mem_la_wdata[2]}),
    .mi({open_n31113,\picorv32_core/pcpi_rs2$26$ }),
    .sr(resetn_placeOpt_12),
    .fx({open_n31117,mem_la_wdata[26]}),
    .q({open_n31118,\uart/uart_bsrr [26]}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*~(B)*~(C)*~(D)*0+A*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B"),
    //.LUTG0("(~(A)*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*~(B)*~(C)*~(D)*1+A*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b0000110000001100),
    .INIT_LUTG0(16'b0111001101100010),
    .INIT_LUTG1(16'b1111110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg2_b8|uart/reg2_b24  (
    .a({open_n31119,\picorv32_core/mem_wordsize [0]}),
    .b({\picorv32_core/pcpi_rs2$8$ ,\picorv32_core/mem_wordsize [1]}),
    .c({\picorv32_core/mem_wordsize [1],mem_la_wdata[0]}),
    .ce(\uart/mux12_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({open_n31120,\picorv32_core/pcpi_rs2$24$ }),
    .e({mem_la_wdata[0],\picorv32_core/pcpi_rs2$8$ }),
    .sr(resetn),
    .f({mem_la_wdata[8],mem_la_wdata[24]}),
    .q({\uart/uart_bsrr [8],\uart/uart_bsrr [24]}));  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)*~(~0*~C))"),
    //.LUTF1("0"),
    //.LUTG0("(~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)*~(~1*~C))"),
    //.LUTG1("D*A*C*~B+D*A*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000001110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0010001001110111),
    .INIT_LUTG1(16'b1010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \uart/reg3_b0|_al_u892  (
    .a({\uart/n9_lutinv ,_al_u700_o}),
    .b({open_n31138,\picorv32_core/pcpi_rs1$3$ }),
    .c({_al_u1179_o,mem_la_addr[2]}),
    .ce(\uart/mux15_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u1175_o,\picorv32_core/n30 [1]}),
    .e({_al_u1168_o,\uart/uart_odr [0]}),
    .mi({mem_la_wdata[0],open_n31140}),
    .f({\uart/mux15_b0_sel_is_2_o ,_al_u892_o}),
    .q({\uart/uart_odr [0],open_n31156}));  // ../src/uart.v(102)
  // ../src/uart.v(102)
  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(~A)"),
    //.LUT1("(~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010101010101),
    .INIT_LUT1(16'b0101010101010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \uart/reg3_b3|uart/reg3_b6  (
    .a({mem_la_wdata[3],mem_la_wdata[6]}),
    .ce(\uart/mux15_b0_sel_is_2_o ),
    .clk(clk_pad),
    .mi({mem_la_wdata[3],mem_la_wdata[6]}),
    .f({n17[3],n17[6]}),
    .q({\uart/uart_odr [3],\uart/uart_odr [6]}));  // ../src/uart.v(102)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*A*~(D*C*~B))"),
    //.LUTF1("(~D)"),
    //.LUTG0("(1*A*~(D*C*~B))"),
    //.LUTG1("(~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b1000101010101010),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \uart/reg3_b5|_al_u1111  (
    .a({open_n31177,_al_u1110_o}),
    .b({open_n31178,\uart/uart_odr [5]}),
    .c({open_n31179,\uart/uart_status_txd [0]}),
    .ce(\uart/mux15_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({mem_la_wdata[5],\uart/uart_status_txd [1]}),
    .e({open_n31180,\uart/uart_status_txd [2]}),
    .mi({mem_la_wdata[5],open_n31182}),
    .f({n17[5],_al_u1111_o}),
    .q({\uart/uart_odr [5],open_n31198}));  // ../src/uart.v(102)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+A*~(B)*C*D*~(0)+A*B*C*~(D)*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+A*B*C*D*0)"),
    //.LUT1("(A*~(B)*D*~(C)*~(1)+~(A)*B*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+A*~(B)*D*C*~(1)+A*B*D*~(C)*1+~(A)*B*~(D)*C*1+A*B*~(D)*C*1+A*B*D*C*1)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010111111100000),
    .INIT_LUT1(16'b1000100011000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg4_b0  (
    .a({\uart/n35 [0],\uart/n35 [0]}),
    .b({_al_u799_o,_al_u799_o}),
    .c({\uart/uart_status_txd [0],_al_u1076_o}),
    .ce(\uart/n30 ),
    .clk(clk_pad),
    .d({_al_u1076_o,\uart/uart_status_txd [0]}),
    .mi({open_n31209,\uart/uart_status_txd [3]}),
    .sr(resetn_placeOpt_1),
    .q({open_n31215,\uart/uart_status_txd [0]}));  // ../src/uart.v(145)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*C*(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B))"),
    //.LUTF1("~C*~B*~D*~A+C*~B*~D*~A+~C*~B*D*~A+C*~B*D*~A+~C*~B*~D*A+C*~B*~D*A+~C*~B*D*A+C*~B*D*A"),
    //.LUTG0("(A*C*(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B))"),
    //.LUTG1("~C*~B*~D*~A+C*~B*~D*~A+C*B*~D*~A+~C*~B*D*~A+C*~B*D*~A+~C*~B*~D*A+C*~B*~D*A+C*B*~D*A+~C*~B*D*A+C*~B*D*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000000000),
    .INIT_LUTF1(16'b0011001100110011),
    .INIT_LUTG0(16'b1010000010000000),
    .INIT_LUTG1(16'b0011001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg4_b1|_al_u893  (
    .a({open_n31216,\uart/n30 }),
    .b({_al_u1081_o,_al_u700_o}),
    .c({_al_u1076_o,mem_la_addr[2]}),
    .ce(\uart/n30 ),
    .clk(clk_pad),
    .d({_al_u1079_o,\picorv32_core/n30 [1]}),
    .e({\uart/n35 [1],\picorv32_core/pcpi_rs1$3$ }),
    .sr(resetn),
    .f({open_n31231,_al_u893_o}),
    .q({\uart/uart_status_txd [1],open_n31235}));  // ../src/uart.v(145)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(A*~(0*D))))"),
    //.LUT1("(B*~(C*~(A*~(1*D))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010001100),
    .INIT_LUT1(16'b0000110010001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg4_b3  (
    .a({\uart/n35 [3],\uart/n35 [3]}),
    .b({_al_u1077_o,_al_u1077_o}),
    .c({_al_u1076_o,_al_u1076_o}),
    .ce(\uart/n30 ),
    .clk(clk_pad),
    .d({\uart/uart_status_txd [1],\uart/uart_status_txd [1]}),
    .mi({open_n31246,\uart/uart_status_txd [3]}),
    .sr(resetn_placeOpt_1),
    .q({open_n31252,\uart/uart_status_txd [3]}));  // ../src/uart.v(145)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0*~((D*B))*~(C)+0*(D*B)*~(C)+~(0)*(D*B)*C+0*(D*B)*C))"),
    //.LUT1("(~A*~(1*~((C*B))*~(D)+1*(C*B)*~(D)+~(1)*(C*B)*D+1*(C*B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010101010101),
    .INIT_LUT1(16'b0001010100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg5_b0  (
    .a({_al_u1164_o,_al_u1164_o}),
    .b({\uart/n51_lutinv ,\uart/n51_lutinv }),
    .c({_al_u1165_o,_al_u1065_o}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({_al_u1065_o,_al_u1165_o}),
    .mi({open_n31263,\uart/uart_status_rxd [3]}),
    .sr(resetn_placeOpt_9),
    .q({open_n31269,\uart/uart_status_rxd [0]}));  // ../src/uart.v(263)
  // ../src/uart.v(263)
  // ../src/uart.v(263)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*(~(A)*~(C)*~(D)*~(0)+A*~(C)*~(D)*~(0)+~(A)*C*~(D)*~(0)+~(A)*~(C)*D*~(0)+A*~(C)*D*~(0)+~(A)*C*D*~(0)+A*C*D*~(0)+~(A)*~(C)*~(D)*0+A*~(C)*~(D)*0+~(A)*C*~(D)*0+A*C*~(D)*0+~(A)*C*D*0))"),
    //.LUTF1("~(~B*D*~(0*C*A))"),
    //.LUTG0("~(~B*(~(A)*~(C)*~(D)*~(1)+A*~(C)*~(D)*~(1)+~(A)*C*~(D)*~(1)+~(A)*~(C)*D*~(1)+A*~(C)*D*~(1)+~(A)*C*D*~(1)+A*C*D*~(1)+~(A)*~(C)*~(D)*1+A*~(C)*~(D)*1+~(A)*C*~(D)*1+A*C*~(D)*1+~(A)*C*D*1))"),
    //.LUTG1("~(~B*D*~(1*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1100110011111111),
    .INIT_LUTG0(16'b1110111111001100),
    .INIT_LUTG1(16'b1110110011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg5_b1|uart/reg5_b3  (
    .a({\uart/mux37_b0_sel_is_3_o ,\uart/n77 [3]}),
    .b({_al_u1160_o,_al_u1160_o}),
    .c({_al_u1070_o,\uart/n51_lutinv }),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({_al_u1189_o,_al_u1065_o}),
    .e({\uart/uart_status_rxd [0],\uart/uart_status_rxd [3]}),
    .sr(resetn_placeOpt_9),
    .q({\uart/uart_status_rxd [1],\uart/uart_status_rxd [3]}));  // ../src/uart.v(263)
  // ../src/uart.v(263)
  // ../src/uart.v(263)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(D)*~((C*B*A))+0*D*~((C*B*A))+~(0)*D*(C*B*A)+0*D*(C*B*A))"),
    //.LUTF1("~(0*~(D)*~((C*~A*B))+0*D*~((C*~A*B))+~(0)*D*(C*~A*B)+0*D*(C*~A*B))"),
    //.LUTG0("~(1*~(D)*~((C*B*A))+1*D*~((C*B*A))+~(1)*D*(C*B*A)+1*D*(C*B*A))"),
    //.LUTG1("~(1*~(D)*~((C*~A*B))+1*D*~((C*~A*B))+~(1)*D*(C*~A*B)+1*D*(C*~A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b1011111111111111),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0000000001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg6_b1|uart/reg6_b3  (
    .a({\uart/n57 [1],_al_u1238_o}),
    .b({_al_u1238_o,\uart/n57 [1]}),
    .c({\uart/n57 [0],\uart/n57 [0]}),
    .ce(\uart/mux51_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({_al_u1086_o,_al_u1086_o}),
    .e({\uart/uart_idr_t [1],\uart/uart_idr_t [3]}),
    .mi({\uart/uart_idr_t [1],\uart/uart_idr_t [3]}),
    .sr(resetn_placeOpt_9),
    .f({_al_u1251_o,_al_u1239_o}),
    .q({\uart/uart_idr [1],\uart/uart_idr [3]}));  // ../src/uart.v(263)
  // ../src/uart.v(263)
  // ../src/uart.v(263)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(D)*~((C*B*A))+0*D*~((C*B*A))+~(0)*D*(C*B*A)+0*D*(C*B*A))"),
    //.LUTF1("~(0*~(C)*~((~D*~B*A))+0*C*~((~D*~B*A))+~(0)*C*(~D*~B*A)+0*C*(~D*~B*A))"),
    //.LUTG0("~(1*~(D)*~((C*B*A))+1*D*~((C*B*A))+~(1)*D*(C*B*A)+1*D*(C*B*A))"),
    //.LUTG1("~(1*~(C)*~((~D*~B*A))+1*C*~((~D*~B*A))+~(1)*C*(~D*~B*A)+1*C*(~D*~B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b1111111111011111),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg6_b4|uart/reg6_b7  (
    .a({_al_u1235_o,_al_u1235_o}),
    .b({\uart/n57 [1],\uart/n57 [1]}),
    .c({_al_u1086_o,\uart/n57 [0]}),
    .ce(\uart/mux51_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\uart/n57 [0],_al_u1086_o}),
    .e({\uart/uart_idr_t [4],\uart/uart_idr_t [7]}),
    .mi({\uart/uart_idr_t [4],\uart/uart_idr_t [7]}),
    .sr(resetn_placeOpt_9),
    .f({_al_u1245_o,_al_u1236_o}),
    .q({\uart/uart_idr [4],\uart/uart_idr [7]}));  // ../src/uart.v(263)
  // ../src/uart.v(263)
  // ../src/uart.v(263)
  EG_PHY_LSLICE #(
    //.LUTF0("~(0*~(D)*~((~C*B*A))+0*D*~((~C*B*A))+~(0)*D*(~C*B*A)+0*D*(~C*B*A))"),
    //.LUTF1("~(0*~(D)*~((C*~A*B))+0*D*~((C*~A*B))+~(0)*D*(C*~A*B)+0*D*(C*~A*B))"),
    //.LUTG0("~(1*~(D)*~((~C*B*A))+1*D*~((~C*B*A))+~(1)*D*(~C*B*A)+1*D*(~C*B*A))"),
    //.LUTG1("~(1*~(D)*~((C*~A*B))+1*D*~((C*~A*B))+~(1)*D*(C*~A*B)+1*D*(C*~A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011111111111),
    .INIT_LUTF1(16'b1011111111111111),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000000001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg6_b5|uart/reg6_b6  (
    .a({\uart/n57 [1],_al_u1235_o}),
    .b({_al_u1235_o,\uart/n57 [1]}),
    .c({\uart/n57 [0],\uart/n57 [0]}),
    .ce(\uart/mux51_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({_al_u1086_o,_al_u1086_o}),
    .e({\uart/uart_idr_t [5],\uart/uart_idr_t [6]}),
    .mi({\uart/uart_idr_t [5],\uart/uart_idr_t [6]}),
    .sr(resetn_placeOpt_9),
    .f({_al_u1249_o,_al_u1241_o}),
    .q({\uart/uart_idr [5],\uart/uart_idr [6]}));  // ../src/uart.v(263)
  // ../src/uart.v(263)
  // ../src/uart.v(263)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+A*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0+A*B*C*D*0)"),
    //.LUTF1("(~(C)*~(A)*~(B)*~(D)*~(0)+~(C)*~(A)*B*~(D)*~(0)+~(C)*A*~(B)*D*~(0)+~(C)*A*B*D*~(0)+~(C)*~(A)*~(B)*~(D)*0+~(C)*~(A)*B*~(D)*0+~(C)*A*B*~(D)*0+C*A*B*~(D)*0+~(C)*~(A)*~(B)*D*0+C*~(A)*~(B)*D*0+~(C)*A*~(B)*D*0+~(C)*~(A)*B*D*0+C*~(A)*B*D*0+~(C)*A*B*D*0+C*A*B*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+A*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1+A*B*C*D*1)"),
    //.LUTG1("(~(C)*~(A)*~(B)*~(D)*~(1)+~(C)*~(A)*B*~(D)*~(1)+~(C)*A*~(B)*D*~(1)+~(C)*A*B*D*~(1)+~(C)*~(A)*~(B)*~(D)*1+~(C)*~(A)*B*~(D)*1+~(C)*A*B*~(D)*1+C*A*B*~(D)*1+~(C)*~(A)*~(B)*D*1+C*~(A)*~(B)*D*1+~(C)*A*~(B)*D*1+~(C)*~(A)*B*D*1+C*~(A)*B*D*1+~(C)*A*B*D*1+C*A*B*D*1)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b0000101000000101),
    .INIT_LUTG0(16'b1111011111010001),
    .INIT_LUTG1(16'b1101111110001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg7_b0|uart/reg7_b5  (
    .a({_al_u1065_o,_al_u1249_o}),
    .b({_al_u1165_o,_al_u1065_o}),
    .c({_al_u1247_o,_al_u1165_o}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({\uart/uart_status_rxd [3],\uart/uart_status_rxd [3]}),
    .e({\uart/uart_idr_t [0],\uart/uart_idr_t [5]}),
    .sr(resetn_placeOpt_9),
    .q({\uart/uart_idr_t [0],\uart/uart_idr_t [5]}));  // ../src/uart.v(263)
  // ../src/uart.v(263)
  // ../src/uart.v(263)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+A*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0+A*B*C*D*0)"),
    //.LUTF1("(~(C)*~(B)*~(A)*~(D)*~(0)+~(C)*~(B)*A*~(D)*~(0)+~(C)*B*~(A)*D*~(0)+~(C)*B*A*D*~(0)+~(C)*~(B)*~(A)*~(D)*0+~(C)*~(B)*A*~(D)*0+~(C)*B*A*~(D)*0+C*B*A*~(D)*0+~(C)*~(B)*~(A)*D*0+C*~(B)*~(A)*D*0+~(C)*B*~(A)*D*0+~(C)*~(B)*A*D*0+C*~(B)*A*D*0+~(C)*B*A*D*0+C*B*A*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+~(A)*B*~(C)*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+A*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1+A*B*C*D*1)"),
    //.LUTG1("(~(C)*~(B)*~(A)*~(D)*~(1)+~(C)*~(B)*A*~(D)*~(1)+~(C)*B*~(A)*D*~(1)+~(C)*B*A*D*~(1)+~(C)*~(B)*~(A)*~(D)*1+~(C)*~(B)*A*~(D)*1+~(C)*B*A*~(D)*1+C*B*A*~(D)*1+~(C)*~(B)*~(A)*D*1+C*~(B)*~(A)*D*1+~(C)*B*~(A)*D*1+~(C)*~(B)*A*D*1+C*~(B)*A*D*1+~(C)*B*A*D*1+C*B*A*D*1)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b0000110000000011),
    .INIT_LUTG0(16'b1111011111010001),
    .INIT_LUTG1(16'b1011111110001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg7_b1|uart/reg7_b4  (
    .a({_al_u1165_o,_al_u1245_o}),
    .b({_al_u1065_o,_al_u1065_o}),
    .c({_al_u1251_o,_al_u1165_o}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({\uart/uart_status_rxd [3],\uart/uart_status_rxd [3]}),
    .e({\uart/uart_idr_t [1],\uart/uart_idr_t [4]}),
    .sr(resetn_placeOpt_9),
    .q({\uart/uart_idr_t [1],\uart/uart_idr_t [4]}));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+A*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0+A*B*C*D*0)"),
    //.LUT1("(~(A)*~(C)*~(D)*~(B)*~(1)+~(A)*~(C)*D*~(B)*~(1)+~(A)*C*~(D)*B*~(1)+~(A)*C*D*B*~(1)+~(A)*~(C)*~(D)*~(B)*1+~(A)*~(C)*D*~(B)*1+~(A)*C*D*~(B)*1+A*C*D*~(B)*1+~(A)*~(C)*~(D)*B*1+A*~(C)*~(D)*B*1+~(A)*C*~(D)*B*1+~(A)*~(C)*D*B*1+A*~(C)*D*B*1+~(A)*C*D*B*1+A*C*D*B*1)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010000010001),
    .INIT_LUT1(16'b1111110101001101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg7_b2  (
    .a({_al_u1243_o,_al_u1243_o}),
    .b({\uart/uart_status_rxd [3],_al_u1065_o}),
    .c({_al_u1065_o,_al_u1165_o}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({_al_u1165_o,\uart/uart_status_rxd [3]}),
    .mi({open_n31382,\uart/uart_idr_t [2]}),
    .sr(resetn_placeOpt_9),
    .q({open_n31388,\uart/uart_idr_t [2]}));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+A*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0+A*B*C*D*0)"),
    //.LUT1("(~(A)*~(C)*~(D)*~(B)*~(1)+~(A)*~(C)*D*~(B)*~(1)+~(A)*C*~(D)*B*~(1)+~(A)*C*D*B*~(1)+~(A)*~(C)*~(D)*~(B)*1+~(A)*~(C)*D*~(B)*1+~(A)*C*D*~(B)*1+A*C*D*~(B)*1+~(A)*~(C)*~(D)*B*1+A*~(C)*~(D)*B*1+~(A)*C*~(D)*B*1+~(A)*~(C)*D*B*1+A*~(C)*D*B*1+~(A)*C*D*B*1+A*C*D*B*1)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010000010001),
    .INIT_LUT1(16'b1111110101001101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg7_b3  (
    .a({_al_u1239_o,_al_u1239_o}),
    .b({\uart/uart_status_rxd [3],_al_u1065_o}),
    .c({_al_u1065_o,_al_u1165_o}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({_al_u1165_o,\uart/uart_status_rxd [3]}),
    .mi({open_n31399,\uart/uart_idr_t [3]}),
    .sr(resetn_placeOpt_9),
    .q({open_n31405,\uart/uart_idr_t [3]}));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+A*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0+A*B*C*D*0)"),
    //.LUT1("(~(A)*~(D)*~(C)*~(B)*~(1)+~(A)*~(D)*C*~(B)*~(1)+~(A)*D*~(C)*B*~(1)+~(A)*D*C*B*~(1)+~(A)*~(D)*~(C)*~(B)*1+~(A)*~(D)*C*~(B)*1+~(A)*D*C*~(B)*1+A*D*C*~(B)*1+~(A)*~(D)*~(C)*B*1+A*~(D)*~(C)*B*1+~(A)*D*~(C)*B*1+~(A)*~(D)*C*B*1+A*~(D)*C*B*1+~(A)*D*C*B*1+A*D*C*B*1)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010000010001),
    .INIT_LUT1(16'b1111010011011101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg7_b6  (
    .a({_al_u1241_o,_al_u1241_o}),
    .b({\uart/uart_status_rxd [3],_al_u1065_o}),
    .c({_al_u1165_o,_al_u1165_o}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({_al_u1065_o,\uart/uart_status_rxd [3]}),
    .mi({open_n31416,\uart/uart_idr_t [6]}),
    .sr(resetn_placeOpt_9),
    .q({open_n31422,\uart/uart_idr_t [6]}));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+~(A)*B*~(C)*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+A*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0+A*B*C*D*0)"),
    //.LUT1("(~(A)*~(D)*~(C)*~(B)*~(1)+~(A)*~(D)*C*~(B)*~(1)+~(A)*D*~(C)*B*~(1)+~(A)*D*C*B*~(1)+~(A)*~(D)*~(C)*~(B)*1+~(A)*~(D)*C*~(B)*1+~(A)*D*C*~(B)*1+A*D*C*~(B)*1+~(A)*~(D)*~(C)*B*1+A*~(D)*~(C)*B*1+~(A)*D*~(C)*B*1+~(A)*~(D)*C*B*1+A*~(D)*C*B*1+~(A)*D*C*B*1+A*D*C*B*1)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010000010001),
    .INIT_LUT1(16'b1111010011011101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg7_b7  (
    .a({_al_u1236_o,_al_u1236_o}),
    .b({\uart/uart_status_rxd [3],_al_u1065_o}),
    .c({_al_u1165_o,_al_u1165_o}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({_al_u1065_o,\uart/uart_status_rxd [3]}),
    .mi({open_n31433,\uart/uart_idr_t [7]}),
    .sr(resetn_placeOpt_9),
    .q({open_n31439,\uart/uart_idr_t [7]}));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A*~(~0*D*~C))"),
    //.LUT1("(~B*~A*~(~1*D*~C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000000010001),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg8_b1  (
    .a({_al_u1071_o,_al_u1071_o}),
    .b({_al_u1072_o,_al_u1072_o}),
    .c({_al_u1068_o,_al_u1068_o}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({\uart/uart_status_rxd [3],\uart/uart_status_rxd [3]}),
    .mi({open_n31450,\uart/uart_cnt_rx [1]}),
    .sr(resetn_placeOpt_9),
    .q({open_n31456,\uart/uart_cnt_rx [1]}));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(0*~(D)*~(B)+0*D*~(B)+~(0)*D*B+0*D*B)))"),
    //.LUT1("(~A*~(C*~(1*~(D)*~(B)+1*D*~(B)+~(1)*D*B+1*D*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010100000101),
    .INIT_LUT1(16'b0101010100010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg8_b2  (
    .a({_al_u1067_o,_al_u1067_o}),
    .b({_al_u1068_o,_al_u1068_o}),
    .c({\uart/uart_status_rxd [3],\uart/uart_status_rxd [3]}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({\uart/uart_cnt_rx [1],\uart/uart_cnt_rx [1]}),
    .mi({open_n31467,\uart/uart_cnt_rx [2]}),
    .sr(resetn_placeOpt_9),
    .q({open_n31473,\uart/uart_cnt_rx [2]}));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)*~(0)+B*C*~(D)*~(0)+B*~(C)*D*~(0)+B*C*D*~(0)+~(B)*C*~(D)*0+B*C*~(D)*0+B*C*D*0))"),
    //.LUT1("(~A*(B*~(C)*~(D)*~(1)+B*C*~(D)*~(1)+B*~(C)*D*~(1)+B*C*D*~(1)+~(B)*C*~(D)*1+B*C*~(D)*1+B*C*D*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010001000100),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg9_b1  (
    .a({_al_u1219_o,_al_u1219_o}),
    .b({\uart/n50 [1],\uart/n50 [1]}),
    .c({_al_u1227_o,_al_u1227_o}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({_al_u1068_o,_al_u1068_o}),
    .mi({open_n31484,\uart/uart_status_rxd [3]}),
    .sr(resetn_placeOpt_9),
    .q({open_n31490,\uart/uart_smp_rx [1]}));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)*~(0)+B*C*~(D)*~(0)+B*~(C)*D*~(0)+B*C*D*~(0)+~(B)*C*~(D)*0+B*C*~(D)*0+B*C*D*0))"),
    //.LUT1("(~A*(B*~(C)*~(D)*~(1)+B*C*~(D)*~(1)+B*~(C)*D*~(1)+B*C*D*~(1)+~(B)*C*~(D)*1+B*C*~(D)*1+B*C*D*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010001000100),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg9_b2  (
    .a({_al_u1219_o,_al_u1219_o}),
    .b({\uart/n50 [2],\uart/n50 [2]}),
    .c({_al_u1224_o,_al_u1224_o}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({_al_u1068_o,_al_u1068_o}),
    .mi({open_n31501,\uart/uart_status_rxd [3]}),
    .sr(resetn_placeOpt_9),
    .q({open_n31507,\uart/uart_smp_rx [2]}));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)*~(0)+B*C*~(D)*~(0)+B*~(C)*D*~(0)+B*C*D*~(0)+~(B)*C*~(D)*0+B*C*~(D)*0+B*C*D*0))"),
    //.LUT1("(~A*(B*~(C)*~(D)*~(1)+B*C*~(D)*~(1)+B*~(C)*D*~(1)+B*C*D*~(1)+~(B)*C*~(D)*1+B*C*~(D)*1+B*C*D*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010001000100),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/reg9_b3  (
    .a({_al_u1219_o,_al_u1219_o}),
    .b({\uart/n50 [3],\uart/n50 [3]}),
    .c({_al_u1221_o,_al_u1221_o}),
    .ce(\uart/uart_op_clock ),
    .clk(clk_pad),
    .d({_al_u1068_o,_al_u1068_o}),
    .mi({open_n31518,\uart/uart_status_rxd [3]}),
    .sr(resetn_placeOpt_9),
    .q({open_n31524,\uart/uart_smp_rx [3]}));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.MACRO("uart/sub1/u0|uart/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \uart/sub1/u0|uart/sub1/ucin  (
    .a({\uart/uart_status_rxd [0],1'b0}),
    .b({1'b0,open_n31525}),
    .f({\uart/n57 [0],open_n31545}),
    .fco(\uart/sub1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/sub1/u0|uart/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \uart/sub1/u2|uart/sub1/u1  (
    .a(\uart/uart_status_rxd [2:1]),
    .b(2'b01),
    .fci(\uart/sub1/c1 ),
    .f(\uart/n57 [2:1]),
    .fco(\uart/sub1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("uart/sub1/u0|uart/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \uart/sub1/ucout|uart/sub1/u3  (
    .a({open_n31572,\uart/uart_status_rxd [3]}),
    .b({open_n31573,1'b0}),
    .fci(\uart/sub1/c3 ),
    .f(\uart/n57 [4:3]));
  EG_PHY_MSLICE #(
    //.MACRO("uart/lt0_0|uart/lt0_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \uart/uart_op_clock_reg|uart/lt0_31  (
    .a({1'b0,\uart/uart_bsrr [31]}),
    .b({1'b1,\uart/uart_counter [31]}),
    .ce(\picorv32_core/n407 ),
    .clk(clk_pad),
    .fci(\uart/lt0_c31 ),
    .f({\uart/n2 ,open_n31613}),
    .q({\uart/uart_op_clock ,open_n31617}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~(~0*D)*~((~C*B))*~(A)+~(~0*D)*(~C*B)*~(A)+~(~(~0*D))*(~C*B)*A+~(~0*D)*(~C*B)*A)"),
    //.LUT1("~(~(~1*D)*~((~C*B))*~(A)+~(~1*D)*(~C*B)*~(A)+~(~(~1*D))*(~C*B)*A+~(~1*D)*(~C*B)*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011110100010),
    .INIT_LUT1(16'b1010001010100010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/uart_status_fe_reg  (
    .a({\uart/mux51_b0_sel_is_3_o ,\uart/mux51_b0_sel_is_3_o }),
    .b({_al_u1086_o,_al_u1086_o}),
    .c({\uart/uart_smp_rx [0],\uart/uart_smp_rx [0]}),
    .clk(clk_pad),
    .d({\uart/uart_status_fe ,\uart/uart_status_fe }),
    .mi({open_n31629,\uart/uart_status_rx_clr }),
    .sr(resetn_placeOpt_14),
    .q({open_n31635,\uart/uart_status_fe }));  // ../src/uart.v(263)
  EG_PHY_MSLICE #(
    //.LUT0("(0*C*B*A*D)"),
    //.LUT1("(1*C*B*A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \uart/uart_status_rx_clr_reg  (
    .a({_al_u1168_o,_al_u1168_o}),
    .b({_al_u1175_o,_al_u1175_o}),
    .c({_al_u1172_o,_al_u1172_o}),
    .clk(clk_pad),
    .d({_al_u1124_o,_al_u1124_o}),
    .mi({open_n31647,\uart/u7_sel_is_3_o }),
    .sr(resetn),
    .q({open_n31653,\uart/uart_status_rx_clr }));  // ../src/uart.v(102)

endmodule 

