// Verilog netlist created by TD v4.3.815
// Wed May  8 18:38:38 2019

`timescale 1ns / 1ps
module sysmem_ml  // al_ip/mem_ml.v(14)
  (
  addra,
  cea,
  clka,
  dia,
  rsta,
  wea,
  doa
  );

  input [9:0] addra;  // al_ip/mem_ml.v(19)
  input cea;  // al_ip/mem_ml.v(21)
  input clka;  // al_ip/mem_ml.v(22)
  input [7:0] dia;  // al_ip/mem_ml.v(18)
  input rsta;  // al_ip/mem_ml.v(23)
  input wea;  // al_ip/mem_ml.v(20)
  output [7:0] doa;  // al_ip/mem_ml.v(16)


  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h440F0007078010DB0F000707081161008BF7C71000804710FE87CE9000011100),
    .INIT_01(256'h8527FE0000972627FEFEFE1727FEFEFE10116150F3C72785C72E8727FC18D680),
    .INIT_02(256'h4037053A3F05C4116185FCFDFEFE07274704C7FDFE00972727FEFCFCFC187161),
    .INIT_03(256'h11615035FE9707FC3DFE9707F7FCFEFE4446FE9342FE5337FC1333FC87DC7101),
    .INIT_04(256'h370F8727403F0FFE370F872785F7FE370F87273FFEFDFCFC18D68044004545C4),
    .INIT_05(256'h3B0585C7FEFE330585F72785F7FE350F872785F7FE3F22FEFDE7FEA8263D0FFD),
    .INIT_06(256'h6F0AB7D687FCFC0727FCFE0747804707FCC30710FEFC00DE80540041272726FE),
    .INIT_07(256'h72726D75000D30312E546E696E2D0A20646F615330612D00476F6972534D5632),
    .INIT_08(256'h00000000000000000000000000000000000000000000003030364E3A003A7330),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_1024x8_sub_000000_000 (
    .addra({addra,3'b111}),
    .cea(cea),
    .clka(clka),
    .dia({open_n68,dia}),
    .rsta(rsta),
    .wea(wea),
    .doa({open_n82,doa}));

endmodule 

