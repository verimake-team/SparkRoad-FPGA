// Verilog netlist created by TD v4.3.815
// Tue May 14 16:18:55 2019

`timescale 1ns / 1ps
module system  // ../src/top.v(3)
  (
  clk,
  resetn_i,
  rxd,
  out_byte,
  out_byte_en,
  trap,
  txd
  );

  input clk;  // ../src/top.v(4)
  input resetn_i;  // ../src/top.v(5)
  input rxd;  // ../src/top.v(14)
  output [7:0] out_byte;  // ../src/top.v(7)
  output out_byte_en;  // ../src/top.v(8)
  output trap;  // ../src/top.v(6)
  output txd;  // ../src/top.v(13)

  wire [1:0] initial_reset;  // ../src/top.v(34)
  wire [31:0] mem_la_addr;  // ../src/top.v(29)
  wire [31:0] mem_la_wdata;  // ../src/top.v(30)
  wire [3:0] mem_la_wstrb;  // ../src/top.v(31)
  wire [31:0] mem_rdata;  // ../src/top.v(23)
  wire [31:0] memory_out;  // ../src/top.v(66)
  wire [7:0] n17;
  wire [1:0] n3;
  wire [31:0] \picorv32_core/alu_add_sub ;  // ../src/picorv32.v(1178)
  wire [31:0] \picorv32_core/alu_out ;  // ../src/picorv32.v(1174)
  wire [31:0] \picorv32_core/alu_out_q ;  // ../src/picorv32.v(1174)
  wire [63:0] \picorv32_core/count_cycle ;  // ../src/picorv32.v(145)
  wire [63:0] \picorv32_core/count_instr ;  // ../src/picorv32.v(145)
  wire [7:0] \picorv32_core/cpu_state ;  // ../src/picorv32.v(1134)
  wire [31:0] \picorv32_core/cpuregs_rs1 ;  // ../src/picorv32.v(1254)
  wire [31:0] \picorv32_core/cpuregs_rs1_z ;  // ../src/picorv32.v(1309)
  wire [31:0] \picorv32_core/cpuregs_rs2 ;  // ../src/picorv32.v(1255)
  wire [31:0] \picorv32_core/cpuregs_rs2_z ;  // ../src/picorv32.v(1310)
  wire [31:0] \picorv32_core/cpuregs_wrdata ;  // ../src/picorv32.v(1252)
  wire [31:0] \picorv32_core/decoded_imm ;  // ../src/picorv32.v(620)
  wire [31:0] \picorv32_core/decoded_imm_uj ;  // ../src/picorv32.v(620)
  wire [4:0] \picorv32_core/decoded_rd ;  // ../src/picorv32.v(619)
  wire [4:0] \picorv32_core/decoded_rs1 ;  // ../src/picorv32.v(619)
  wire [4:0] \picorv32_core/decoded_rs2 ;  // ../src/picorv32.v(619)
  wire [4:0] \picorv32_core/latched_rd ;  // ../src/picorv32.v(1163)
  wire [15:0] \picorv32_core/mem_16bit_buffer ;  // ../src/picorv32.v(331)
  wire [31:0] \picorv32_core/mem_rdata_latched ;  // ../src/picorv32.v(334)
  wire [31:0] \picorv32_core/mem_rdata_latched_noshuffle ;  // ../src/picorv32.v(333)
  wire [31:0] \picorv32_core/mem_rdata_q ;  // ../src/picorv32.v(319)
  wire [31:0] \picorv32_core/mem_rdata_word ;  // ../src/picorv32.v(318)
  wire [1:0] \picorv32_core/mem_state ;  // ../src/picorv32.v(316)
  wire [1:0] \picorv32_core/mem_wordsize ;  // ../src/picorv32.v(317)
  wire [4:0] \picorv32_core/n102 ;
  wire [1:0] \picorv32_core/n103 ;
  wire [2:0] \picorv32_core/n105 ;
  wire [4:0] \picorv32_core/n107 ;
  wire [4:0] \picorv32_core/n108 ;
  wire [24:0] \picorv32_core/n109 ;
  wire [24:0] \picorv32_core/n110 ;
  wire [1:0] \picorv32_core/n112 ;
  wire [3:0] \picorv32_core/n116 ;
  wire [1:0] \picorv32_core/n124 ;
  wire [1:0] \picorv32_core/n127 ;
  wire [15:0] \picorv32_core/n128 ;
  wire [15:0] \picorv32_core/n133 ;
  wire [1:0] \picorv32_core/n135 ;
  wire [15:0] \picorv32_core/n136 ;
  wire [1:0] \picorv32_core/n143 ;
  wire [1:0] \picorv32_core/n145 ;
  wire [1:0] \picorv32_core/n146 ;
  wire [1:0] \picorv32_core/n147 ;
  wire [1:0] \picorv32_core/n154 ;
  wire [1:0] \picorv32_core/n186 ;
  wire [2:0] \picorv32_core/n189 ;
  wire [2:0] \picorv32_core/n192 ;
  wire [4:0] \picorv32_core/n195 ;
  wire [4:0] \picorv32_core/n200 ;
  wire [3:0] \picorv32_core/n205 ;
  wire [4:0] \picorv32_core/n206 ;
  wire [4:0] \picorv32_core/n208 ;
  wire [4:0] \picorv32_core/n209 ;
  wire [4:0] \picorv32_core/n212 ;
  wire [4:0] \picorv32_core/n218 ;
  wire [4:0] \picorv32_core/n222 ;
  wire [4:0] \picorv32_core/n225 ;
  wire [4:0] \picorv32_core/n226 ;
  wire [4:0] \picorv32_core/n227 ;
  wire [4:0] \picorv32_core/n229 ;
  wire [4:0] \picorv32_core/n230 ;
  wire [4:0] \picorv32_core/n231 ;
  wire [4:0] \picorv32_core/n235 ;
  wire [4:0] \picorv32_core/n236 ;
  wire [4:0] \picorv32_core/n237 ;
  wire [4:0] \picorv32_core/n245 ;
  wire [4:0] \picorv32_core/n246 ;
  wire [4:0] \picorv32_core/n247 ;
  wire [29:0] \picorv32_core/n248 ;
  wire [29:0] \picorv32_core/n30 ;
  wire [31:0] \picorv32_core/n31 ;
  wire [31:0] \picorv32_core/n32 ;
  wire [31:0] \picorv32_core/n358 ;
  wire [3:0] \picorv32_core/n38 ;
  wire [31:0] \picorv32_core/n39 ;
  wire [3:0] \picorv32_core/n40 ;
  wire [31:0] \picorv32_core/n41 ;
  wire [31:0] \picorv32_core/n42 ;
  wire [31:0] \picorv32_core/n433 ;
  wire [31:0] \picorv32_core/n434 ;
  wire [31:0] \picorv32_core/n439 ;
  wire [31:0] \picorv32_core/n441 ;
  wire [31:0] \picorv32_core/n443 ;
  wire [2:0] \picorv32_core/n449 ;
  wire [4:0] \picorv32_core/n45 ;
  wire [31:0] \picorv32_core/n450 ;
  wire [31:0] \picorv32_core/n453 ;
  wire [31:0] \picorv32_core/n455 ;
  wire [63:0] \picorv32_core/n459 ;
  wire [4:0] \picorv32_core/n47 ;
  wire [3:0] \picorv32_core/n49 ;
  wire [31:0] \picorv32_core/n500 ;
  wire [2:0] \picorv32_core/n501 ;
  wire [31:0] \picorv32_core/n502 ;
  wire [63:0] \picorv32_core/n503 ;
  wire [31:0] \picorv32_core/n504 ;
  wire [31:0] \picorv32_core/n508 ;
  wire [31:0] \picorv32_core/n511 ;
  wire [7:0] \picorv32_core/n516 ;
  wire [31:0] \picorv32_core/n518 ;
  wire [4:0] \picorv32_core/n52 ;
  wire [7:0] \picorv32_core/n521 ;
  wire [7:0] \picorv32_core/n524 ;
  wire [31:0] \picorv32_core/n525 ;
  wire [31:0] \picorv32_core/n527 ;
  wire [31:0] \picorv32_core/n528 ;
  wire [16:0] \picorv32_core/n53 ;
  wire [4:0] \picorv32_core/n532 ;
  wire [31:0] \picorv32_core/n543 ;
  wire [4:0] \picorv32_core/n546 ;
  wire [7:0] \picorv32_core/n549 ;
  wire [9:0] \picorv32_core/n55 ;
  wire [31:0] \picorv32_core/n558 ;
  wire [5:0] \picorv32_core/n559 ;
  wire [31:0] \picorv32_core/n563 ;
  wire [5:0] \picorv32_core/n564 ;
  wire [31:0] \picorv32_core/n565 ;
  wire [4:0] \picorv32_core/n566 ;
  wire [31:0] \picorv32_core/n567 ;
  wire [7:0] \picorv32_core/n569 ;
  wire [9:0] \picorv32_core/n57 ;
  wire [31:0] \picorv32_core/n570 ;
  wire [4:0] \picorv32_core/n571 ;
  wire [1:0] \picorv32_core/n575 ;
  wire [31:0] \picorv32_core/n576 ;
  wire [1:0] \picorv32_core/n583 ;
  wire [31:0] \picorv32_core/n584 ;
  wire [9:0] \picorv32_core/n59 ;
  wire [4:0] \picorv32_core/n60 ;
  wire [1:0] \picorv32_core/n601 ;
  wire [2:0] \picorv32_core/n62 ;
  wire [2:0] \picorv32_core/n64 ;
  wire [31:0] \picorv32_core/n641 ;
  wire [31:0] \picorv32_core/n642 ;
  wire [1:0] \picorv32_core/n652 ;
  wire [31:0] \picorv32_core/n656 ;
  wire [31:0] \picorv32_core/n658 ;
  wire [2:0] \picorv32_core/n66 ;
  wire [7:0] \picorv32_core/n661 ;
  wire [1:0] \picorv32_core/n672 ;
  wire [2:0] \picorv32_core/n68 ;
  wire [4:0] \picorv32_core/n688 ;
  wire [9:0] \picorv32_core/n69 ;
  wire [7:0] \picorv32_core/n692 ;
  wire [31:0] \picorv32_core/n693 ;
  wire [31:0] \picorv32_core/n694 ;
  wire [31:0] \picorv32_core/n695 ;
  wire [4:0] \picorv32_core/n696 ;
  wire [19:0] \picorv32_core/n70 ;
  wire [4:0] \picorv32_core/n71 ;
  wire [7:0] \picorv32_core/n716 ;
  wire [31:0] \picorv32_core/n725 ;
  wire [4:0] \picorv32_core/n726 ;
  wire [4:0] \picorv32_core/n91 ;
  wire [4:0] \picorv32_core/n93 ;
  wire [1:0] \picorv32_core/n94 ;
  wire [2:0] \picorv32_core/n95 ;
  wire [31:0] \picorv32_core/next_pc ;  // ../src/picorv32.v(168)
  wire [31:0] \picorv32_core/reg_next_pc ;  // ../src/picorv32.v(146)
  wire [31:0] \picorv32_core/reg_out ;  // ../src/picorv32.v(146)
  wire [31:0] \picorv32_core/reg_pc ;  // ../src/picorv32.v(146)
  wire [4:0] \picorv32_core/reg_sh ;  // ../src/picorv32.v(151)
  wire  \picorv32_core/sel0_b28/B0 ;
  wire  \picorv32_core/sel0_b28/B2 ;
  wire  \picorv32_core/sel0_b29/B2 ;
  wire  \picorv32_core/sel0_b30/B2 ;
  wire  \picorv32_core/sel0_b31/B2 ;
  wire  \picorv32_core/sel0_b63/B2 ;
  wire  \picorv32_core/sel11_b0/B1 ;
  wire  \picorv32_core/sel11_b0/B3 ;
  wire  \picorv32_core/sel11_b1/B1 ;
  wire  \picorv32_core/sel11_b1/B2 ;
  wire  \picorv32_core/sel11_b1/B3 ;
  wire  \picorv32_core/sel11_b1/B5 ;
  wire  \picorv32_core/sel11_b10/B1 ;
  wire  \picorv32_core/sel11_b10/B2 ;
  wire  \picorv32_core/sel11_b10/B3 ;
  wire  \picorv32_core/sel11_b10/B5 ;
  wire  \picorv32_core/sel11_b11/B1 ;
  wire  \picorv32_core/sel11_b11/B2 ;
  wire  \picorv32_core/sel11_b11/B3 ;
  wire  \picorv32_core/sel11_b11/B5 ;
  wire  \picorv32_core/sel11_b12/B2 ;
  wire  \picorv32_core/sel11_b12/B4 ;
  wire  \picorv32_core/sel11_b12/B5 ;
  wire  \picorv32_core/sel11_b13/B4 ;
  wire  \picorv32_core/sel11_b13/B5 ;
  wire  \picorv32_core/sel11_b14/B4 ;
  wire  \picorv32_core/sel11_b14/B5 ;
  wire  \picorv32_core/sel11_b15/B4 ;
  wire  \picorv32_core/sel11_b15/B5 ;
  wire  \picorv32_core/sel11_b16/B4 ;
  wire  \picorv32_core/sel11_b16/B5 ;
  wire  \picorv32_core/sel11_b17/B4 ;
  wire  \picorv32_core/sel11_b17/B5 ;
  wire  \picorv32_core/sel11_b18/B4 ;
  wire  \picorv32_core/sel11_b18/B5 ;
  wire  \picorv32_core/sel11_b19/B4 ;
  wire  \picorv32_core/sel11_b19/B5 ;
  wire  \picorv32_core/sel11_b2/B1 ;
  wire  \picorv32_core/sel11_b2/B2 ;
  wire  \picorv32_core/sel11_b2/B3 ;
  wire  \picorv32_core/sel11_b2/B5 ;
  wire  \picorv32_core/sel11_b20/B4 ;
  wire  \picorv32_core/sel11_b20/B5 ;
  wire  \picorv32_core/sel11_b21/B4 ;
  wire  \picorv32_core/sel11_b22/B4 ;
  wire  \picorv32_core/sel11_b23/B4 ;
  wire  \picorv32_core/sel11_b24/B4 ;
  wire  \picorv32_core/sel11_b25/B4 ;
  wire  \picorv32_core/sel11_b26/B4 ;
  wire  \picorv32_core/sel11_b27/B4 ;
  wire  \picorv32_core/sel11_b28/B4 ;
  wire  \picorv32_core/sel11_b29/B4 ;
  wire  \picorv32_core/sel11_b3/B1 ;
  wire  \picorv32_core/sel11_b3/B2 ;
  wire  \picorv32_core/sel11_b3/B3 ;
  wire  \picorv32_core/sel11_b3/B5 ;
  wire  \picorv32_core/sel11_b30/B4 ;
  wire  \picorv32_core/sel11_b31/B4 ;
  wire  \picorv32_core/sel11_b4/B1 ;
  wire  \picorv32_core/sel11_b4/B2 ;
  wire  \picorv32_core/sel11_b4/B3 ;
  wire  \picorv32_core/sel11_b4/B5 ;
  wire  \picorv32_core/sel11_b5/B1 ;
  wire  \picorv32_core/sel11_b5/B2 ;
  wire  \picorv32_core/sel11_b5/B3 ;
  wire  \picorv32_core/sel11_b5/B5 ;
  wire  \picorv32_core/sel11_b6/B1 ;
  wire  \picorv32_core/sel11_b6/B2 ;
  wire  \picorv32_core/sel11_b6/B3 ;
  wire  \picorv32_core/sel11_b6/B5 ;
  wire  \picorv32_core/sel11_b7/B1 ;
  wire  \picorv32_core/sel11_b7/B2 ;
  wire  \picorv32_core/sel11_b7/B3 ;
  wire  \picorv32_core/sel11_b7/B5 ;
  wire  \picorv32_core/sel11_b8/B1 ;
  wire  \picorv32_core/sel11_b8/B2 ;
  wire  \picorv32_core/sel11_b8/B3 ;
  wire  \picorv32_core/sel11_b8/B5 ;
  wire  \picorv32_core/sel11_b9/B1 ;
  wire  \picorv32_core/sel11_b9/B2 ;
  wire  \picorv32_core/sel11_b9/B3 ;
  wire  \picorv32_core/sel11_b9/B5 ;
  wire  \picorv32_core/sel12/B0 ;
  wire  \picorv32_core/sel12/B1 ;
  wire  \picorv32_core/sel12/B2 ;
  wire  \picorv32_core/sel12/B3 ;
  wire  \picorv32_core/sel13_b0/B0 ;
  wire  \picorv32_core/sel13_b0/B1 ;
  wire  \picorv32_core/sel13_b0/B2 ;
  wire  \picorv32_core/sel13_b0/B3 ;
  wire  \picorv32_core/sel13_b0/B4 ;
  wire  \picorv32_core/sel13_b1/B0 ;
  wire  \picorv32_core/sel13_b1/B1 ;
  wire  \picorv32_core/sel13_b1/B2 ;
  wire  \picorv32_core/sel13_b1/B4 ;
  wire  \picorv32_core/sel13_b10/B0 ;
  wire  \picorv32_core/sel13_b10/B1 ;
  wire  \picorv32_core/sel13_b10/B2 ;
  wire  \picorv32_core/sel13_b10/B4 ;
  wire  \picorv32_core/sel13_b11/B0 ;
  wire  \picorv32_core/sel13_b11/B1 ;
  wire  \picorv32_core/sel13_b11/B2 ;
  wire  \picorv32_core/sel13_b11/B4 ;
  wire  \picorv32_core/sel13_b12/B0 ;
  wire  \picorv32_core/sel13_b12/B1 ;
  wire  \picorv32_core/sel13_b12/B2 ;
  wire  \picorv32_core/sel13_b12/B4 ;
  wire  \picorv32_core/sel13_b13/B0 ;
  wire  \picorv32_core/sel13_b13/B1 ;
  wire  \picorv32_core/sel13_b13/B2 ;
  wire  \picorv32_core/sel13_b13/B4 ;
  wire  \picorv32_core/sel13_b14/B0 ;
  wire  \picorv32_core/sel13_b14/B1 ;
  wire  \picorv32_core/sel13_b14/B2 ;
  wire  \picorv32_core/sel13_b14/B4 ;
  wire  \picorv32_core/sel13_b15/B0 ;
  wire  \picorv32_core/sel13_b15/B1 ;
  wire  \picorv32_core/sel13_b15/B2 ;
  wire  \picorv32_core/sel13_b15/B4 ;
  wire  \picorv32_core/sel13_b16/B0 ;
  wire  \picorv32_core/sel13_b16/B1 ;
  wire  \picorv32_core/sel13_b16/B2 ;
  wire  \picorv32_core/sel13_b16/B4 ;
  wire  \picorv32_core/sel13_b17/B0 ;
  wire  \picorv32_core/sel13_b17/B1 ;
  wire  \picorv32_core/sel13_b17/B2 ;
  wire  \picorv32_core/sel13_b17/B4 ;
  wire  \picorv32_core/sel13_b18/B0 ;
  wire  \picorv32_core/sel13_b18/B1 ;
  wire  \picorv32_core/sel13_b18/B2 ;
  wire  \picorv32_core/sel13_b18/B4 ;
  wire  \picorv32_core/sel13_b19/B0 ;
  wire  \picorv32_core/sel13_b19/B1 ;
  wire  \picorv32_core/sel13_b19/B2 ;
  wire  \picorv32_core/sel13_b19/B4 ;
  wire  \picorv32_core/sel13_b2/B0 ;
  wire  \picorv32_core/sel13_b2/B1 ;
  wire  \picorv32_core/sel13_b2/B2 ;
  wire  \picorv32_core/sel13_b2/B4 ;
  wire  \picorv32_core/sel13_b20/B0 ;
  wire  \picorv32_core/sel13_b20/B1 ;
  wire  \picorv32_core/sel13_b20/B2 ;
  wire  \picorv32_core/sel13_b20/B4 ;
  wire  \picorv32_core/sel13_b21/B0 ;
  wire  \picorv32_core/sel13_b21/B1 ;
  wire  \picorv32_core/sel13_b21/B2 ;
  wire  \picorv32_core/sel13_b21/B4 ;
  wire  \picorv32_core/sel13_b22/B0 ;
  wire  \picorv32_core/sel13_b22/B1 ;
  wire  \picorv32_core/sel13_b22/B2 ;
  wire  \picorv32_core/sel13_b22/B4 ;
  wire  \picorv32_core/sel13_b23/B0 ;
  wire  \picorv32_core/sel13_b23/B1 ;
  wire  \picorv32_core/sel13_b23/B2 ;
  wire  \picorv32_core/sel13_b23/B4 ;
  wire  \picorv32_core/sel13_b24/B0 ;
  wire  \picorv32_core/sel13_b24/B1 ;
  wire  \picorv32_core/sel13_b24/B2 ;
  wire  \picorv32_core/sel13_b24/B4 ;
  wire  \picorv32_core/sel13_b25/B0 ;
  wire  \picorv32_core/sel13_b25/B1 ;
  wire  \picorv32_core/sel13_b25/B2 ;
  wire  \picorv32_core/sel13_b25/B4 ;
  wire  \picorv32_core/sel13_b26/B0 ;
  wire  \picorv32_core/sel13_b26/B1 ;
  wire  \picorv32_core/sel13_b26/B2 ;
  wire  \picorv32_core/sel13_b26/B4 ;
  wire  \picorv32_core/sel13_b27/B0 ;
  wire  \picorv32_core/sel13_b27/B1 ;
  wire  \picorv32_core/sel13_b27/B2 ;
  wire  \picorv32_core/sel13_b27/B4 ;
  wire  \picorv32_core/sel13_b28/B0 ;
  wire  \picorv32_core/sel13_b28/B1 ;
  wire  \picorv32_core/sel13_b28/B2 ;
  wire  \picorv32_core/sel13_b28/B4 ;
  wire  \picorv32_core/sel13_b29/B0 ;
  wire  \picorv32_core/sel13_b29/B1 ;
  wire  \picorv32_core/sel13_b29/B2 ;
  wire  \picorv32_core/sel13_b29/B4 ;
  wire  \picorv32_core/sel13_b3/B0 ;
  wire  \picorv32_core/sel13_b3/B1 ;
  wire  \picorv32_core/sel13_b3/B2 ;
  wire  \picorv32_core/sel13_b3/B4 ;
  wire  \picorv32_core/sel13_b30/B0 ;
  wire  \picorv32_core/sel13_b30/B1 ;
  wire  \picorv32_core/sel13_b30/B2 ;
  wire  \picorv32_core/sel13_b30/B4 ;
  wire  \picorv32_core/sel13_b31/B0 ;
  wire  \picorv32_core/sel13_b31/B1 ;
  wire  \picorv32_core/sel13_b31/B2 ;
  wire  \picorv32_core/sel13_b31/B4 ;
  wire  \picorv32_core/sel13_b4/B0 ;
  wire  \picorv32_core/sel13_b4/B1 ;
  wire  \picorv32_core/sel13_b4/B2 ;
  wire  \picorv32_core/sel13_b4/B4 ;
  wire  \picorv32_core/sel13_b5/B0 ;
  wire  \picorv32_core/sel13_b5/B1 ;
  wire  \picorv32_core/sel13_b5/B2 ;
  wire  \picorv32_core/sel13_b5/B4 ;
  wire  \picorv32_core/sel13_b6/B0 ;
  wire  \picorv32_core/sel13_b6/B1 ;
  wire  \picorv32_core/sel13_b6/B2 ;
  wire  \picorv32_core/sel13_b6/B4 ;
  wire  \picorv32_core/sel13_b7/B0 ;
  wire  \picorv32_core/sel13_b7/B1 ;
  wire  \picorv32_core/sel13_b7/B2 ;
  wire  \picorv32_core/sel13_b7/B4 ;
  wire  \picorv32_core/sel13_b8/B0 ;
  wire  \picorv32_core/sel13_b8/B1 ;
  wire  \picorv32_core/sel13_b8/B2 ;
  wire  \picorv32_core/sel13_b8/B4 ;
  wire  \picorv32_core/sel13_b9/B0 ;
  wire  \picorv32_core/sel13_b9/B1 ;
  wire  \picorv32_core/sel13_b9/B2 ;
  wire  \picorv32_core/sel13_b9/B4 ;
  wire  \picorv32_core/sel16_b0/B0 ;
  wire  \picorv32_core/sel16_b0/B1 ;
  wire  \picorv32_core/sel16_b0/B2 ;
  wire  \picorv32_core/sel16_b0/B3 ;
  wire  \picorv32_core/sel16_b1/B0 ;
  wire  \picorv32_core/sel16_b1/B1 ;
  wire  \picorv32_core/sel16_b1/B2 ;
  wire  \picorv32_core/sel16_b1/B3 ;
  wire  \picorv32_core/sel16_b10/B0 ;
  wire  \picorv32_core/sel16_b10/B1 ;
  wire  \picorv32_core/sel16_b10/B2 ;
  wire  \picorv32_core/sel16_b10/B3 ;
  wire  \picorv32_core/sel16_b11/B0 ;
  wire  \picorv32_core/sel16_b11/B1 ;
  wire  \picorv32_core/sel16_b11/B2 ;
  wire  \picorv32_core/sel16_b11/B3 ;
  wire  \picorv32_core/sel16_b12/B0 ;
  wire  \picorv32_core/sel16_b12/B1 ;
  wire  \picorv32_core/sel16_b12/B2 ;
  wire  \picorv32_core/sel16_b12/B3 ;
  wire  \picorv32_core/sel16_b13/B0 ;
  wire  \picorv32_core/sel16_b13/B1 ;
  wire  \picorv32_core/sel16_b13/B2 ;
  wire  \picorv32_core/sel16_b13/B3 ;
  wire  \picorv32_core/sel16_b14/B0 ;
  wire  \picorv32_core/sel16_b14/B1 ;
  wire  \picorv32_core/sel16_b14/B2 ;
  wire  \picorv32_core/sel16_b14/B3 ;
  wire  \picorv32_core/sel16_b15/B0 ;
  wire  \picorv32_core/sel16_b15/B1 ;
  wire  \picorv32_core/sel16_b15/B2 ;
  wire  \picorv32_core/sel16_b15/B3 ;
  wire  \picorv32_core/sel16_b16/B0 ;
  wire  \picorv32_core/sel16_b16/B1 ;
  wire  \picorv32_core/sel16_b16/B2 ;
  wire  \picorv32_core/sel16_b16/B3 ;
  wire  \picorv32_core/sel16_b17/B0 ;
  wire  \picorv32_core/sel16_b17/B1 ;
  wire  \picorv32_core/sel16_b17/B2 ;
  wire  \picorv32_core/sel16_b17/B3 ;
  wire  \picorv32_core/sel16_b18/B0 ;
  wire  \picorv32_core/sel16_b18/B1 ;
  wire  \picorv32_core/sel16_b18/B2 ;
  wire  \picorv32_core/sel16_b18/B3 ;
  wire  \picorv32_core/sel16_b19/B0 ;
  wire  \picorv32_core/sel16_b19/B1 ;
  wire  \picorv32_core/sel16_b19/B2 ;
  wire  \picorv32_core/sel16_b19/B3 ;
  wire  \picorv32_core/sel16_b2/B0 ;
  wire  \picorv32_core/sel16_b2/B1 ;
  wire  \picorv32_core/sel16_b2/B2 ;
  wire  \picorv32_core/sel16_b2/B3 ;
  wire  \picorv32_core/sel16_b20/B0 ;
  wire  \picorv32_core/sel16_b20/B1 ;
  wire  \picorv32_core/sel16_b20/B2 ;
  wire  \picorv32_core/sel16_b20/B3 ;
  wire  \picorv32_core/sel16_b21/B0 ;
  wire  \picorv32_core/sel16_b21/B1 ;
  wire  \picorv32_core/sel16_b21/B2 ;
  wire  \picorv32_core/sel16_b21/B3 ;
  wire  \picorv32_core/sel16_b22/B0 ;
  wire  \picorv32_core/sel16_b22/B1 ;
  wire  \picorv32_core/sel16_b22/B2 ;
  wire  \picorv32_core/sel16_b22/B3 ;
  wire  \picorv32_core/sel16_b23/B0 ;
  wire  \picorv32_core/sel16_b23/B1 ;
  wire  \picorv32_core/sel16_b23/B2 ;
  wire  \picorv32_core/sel16_b23/B3 ;
  wire  \picorv32_core/sel16_b24/B0 ;
  wire  \picorv32_core/sel16_b24/B1 ;
  wire  \picorv32_core/sel16_b24/B2 ;
  wire  \picorv32_core/sel16_b24/B3 ;
  wire  \picorv32_core/sel16_b25/B0 ;
  wire  \picorv32_core/sel16_b25/B1 ;
  wire  \picorv32_core/sel16_b25/B2 ;
  wire  \picorv32_core/sel16_b25/B3 ;
  wire  \picorv32_core/sel16_b26/B0 ;
  wire  \picorv32_core/sel16_b26/B1 ;
  wire  \picorv32_core/sel16_b26/B2 ;
  wire  \picorv32_core/sel16_b26/B3 ;
  wire  \picorv32_core/sel16_b27/B0 ;
  wire  \picorv32_core/sel16_b27/B1 ;
  wire  \picorv32_core/sel16_b27/B2 ;
  wire  \picorv32_core/sel16_b27/B3 ;
  wire  \picorv32_core/sel16_b28/B0 ;
  wire  \picorv32_core/sel16_b28/B1 ;
  wire  \picorv32_core/sel16_b28/B2 ;
  wire  \picorv32_core/sel16_b28/B3 ;
  wire  \picorv32_core/sel16_b29/B0 ;
  wire  \picorv32_core/sel16_b29/B1 ;
  wire  \picorv32_core/sel16_b29/B2 ;
  wire  \picorv32_core/sel16_b29/B3 ;
  wire  \picorv32_core/sel16_b3/B0 ;
  wire  \picorv32_core/sel16_b3/B1 ;
  wire  \picorv32_core/sel16_b3/B2 ;
  wire  \picorv32_core/sel16_b3/B3 ;
  wire  \picorv32_core/sel16_b30/B0 ;
  wire  \picorv32_core/sel16_b30/B1 ;
  wire  \picorv32_core/sel16_b30/B2 ;
  wire  \picorv32_core/sel16_b30/B3 ;
  wire  \picorv32_core/sel16_b31/B0 ;
  wire  \picorv32_core/sel16_b31/B1 ;
  wire  \picorv32_core/sel16_b31/B2 ;
  wire  \picorv32_core/sel16_b31/B3 ;
  wire  \picorv32_core/sel16_b4/B0 ;
  wire  \picorv32_core/sel16_b4/B1 ;
  wire  \picorv32_core/sel16_b4/B2 ;
  wire  \picorv32_core/sel16_b4/B3 ;
  wire  \picorv32_core/sel16_b5/B0 ;
  wire  \picorv32_core/sel16_b5/B1 ;
  wire  \picorv32_core/sel16_b5/B2 ;
  wire  \picorv32_core/sel16_b5/B3 ;
  wire  \picorv32_core/sel16_b6/B0 ;
  wire  \picorv32_core/sel16_b6/B1 ;
  wire  \picorv32_core/sel16_b6/B2 ;
  wire  \picorv32_core/sel16_b6/B3 ;
  wire  \picorv32_core/sel16_b7/B0 ;
  wire  \picorv32_core/sel16_b7/B1 ;
  wire  \picorv32_core/sel16_b7/B2 ;
  wire  \picorv32_core/sel16_b7/B3 ;
  wire  \picorv32_core/sel16_b8/B0 ;
  wire  \picorv32_core/sel16_b8/B1 ;
  wire  \picorv32_core/sel16_b8/B2 ;
  wire  \picorv32_core/sel16_b8/B3 ;
  wire  \picorv32_core/sel16_b9/B0 ;
  wire  \picorv32_core/sel16_b9/B1 ;
  wire  \picorv32_core/sel16_b9/B2 ;
  wire  \picorv32_core/sel16_b9/B3 ;
  wire  \picorv32_core/sel18/B0 ;
  wire  \picorv32_core/sel18/B1 ;
  wire  \picorv32_core/sel19_b2/B0 ;
  wire  \picorv32_core/sel19_b3/B0 ;
  wire  \picorv32_core/sel1_b0/B0 ;
  wire  \picorv32_core/sel1_b0/B1 ;
  wire  \picorv32_core/sel1_b1/B0 ;
  wire  \picorv32_core/sel1_b1/B1 ;
  wire  \picorv32_core/sel1_b2/B0 ;
  wire  \picorv32_core/sel1_b2/B1 ;
  wire  \picorv32_core/sel1_b3/B0 ;
  wire  \picorv32_core/sel1_b3/B1 ;
  wire  \picorv32_core/sel1_b4/B0 ;
  wire  \picorv32_core/sel1_b4/B1 ;
  wire  \picorv32_core/sel2/B0 ;
  wire  \picorv32_core/sel2/B1 ;
  wire  \picorv32_core/sel2/B2 ;
  wire  \picorv32_core/sel23/B0 ;
  wire  \picorv32_core/sel23/B2 ;
  wire  \picorv32_core/sel23/B3 ;
  wire  \picorv32_core/sel27_b16/B0 ;
  wire  \picorv32_core/sel27_b16/B1 ;
  wire  \picorv32_core/sel27_b16/B2 ;
  wire  \picorv32_core/sel27_b17/B2 ;
  wire  \picorv32_core/sel27_b18/B2 ;
  wire  \picorv32_core/sel27_b19/B2 ;
  wire  \picorv32_core/sel27_b20/B2 ;
  wire  \picorv32_core/sel27_b21/B2 ;
  wire  \picorv32_core/sel27_b22/B2 ;
  wire  \picorv32_core/sel27_b23/B2 ;
  wire  \picorv32_core/sel27_b24/B2 ;
  wire  \picorv32_core/sel27_b25/B2 ;
  wire  \picorv32_core/sel27_b26/B2 ;
  wire  \picorv32_core/sel27_b27/B2 ;
  wire  \picorv32_core/sel27_b28/B2 ;
  wire  \picorv32_core/sel27_b29/B2 ;
  wire  \picorv32_core/sel27_b30/B2 ;
  wire  \picorv32_core/sel27_b31/B2 ;
  wire  \picorv32_core/sel28/B0 ;
  wire  \picorv32_core/sel28/B1 ;
  wire  \picorv32_core/sel28/B2 ;
  wire  \picorv32_core/sel28/B3 ;
  wire  \picorv32_core/sel28/B4 ;
  wire  \picorv32_core/sel29_b0/B0 ;
  wire  \picorv32_core/sel29_b0/B1 ;
  wire  \picorv32_core/sel29_b0/B2 ;
  wire  \picorv32_core/sel29_b0/B3 ;
  wire  \picorv32_core/sel29_b0/B4 ;
  wire  \picorv32_core/sel29_b0/B5 ;
  wire  \picorv32_core/sel29_b0/B7 ;
  wire  \picorv32_core/sel29_b1/B0 ;
  wire  \picorv32_core/sel29_b1/B1 ;
  wire  \picorv32_core/sel29_b1/B2 ;
  wire  \picorv32_core/sel29_b1/B3 ;
  wire  \picorv32_core/sel29_b1/B4 ;
  wire  \picorv32_core/sel29_b1/B5 ;
  wire  \picorv32_core/sel29_b1/B7 ;
  wire  \picorv32_core/sel32/B1 ;
  wire  \picorv32_core/sel32/B2 ;
  wire  \picorv32_core/sel32/B4 ;
  wire  \picorv32_core/sel33/B0 ;
  wire  \picorv32_core/sel33/B2 ;
  wire  \picorv32_core/sel34/B0 ;
  wire  \picorv32_core/sel34/B1 ;
  wire  \picorv32_core/sel34/B2 ;
  wire  \picorv32_core/sel35/B0 ;
  wire  \picorv32_core/sel35/B2 ;
  wire  \picorv32_core/sel36/B0 ;
  wire  \picorv32_core/sel36/B2 ;
  wire  \picorv32_core/sel37/B0 ;
  wire  \picorv32_core/sel37/B2 ;
  wire  \picorv32_core/sel38_b0/B0 ;
  wire  \picorv32_core/sel38_b0/B1 ;
  wire  \picorv32_core/sel38_b0/B2 ;
  wire  \picorv32_core/sel38_b0/B3 ;
  wire  \picorv32_core/sel38_b0/B4 ;
  wire  \picorv32_core/sel38_b0/B5 ;
  wire  \picorv32_core/sel38_b0/B6 ;
  wire  \picorv32_core/sel38_b0/B7 ;
  wire  \picorv32_core/sel38_b1/B0 ;
  wire  \picorv32_core/sel38_b1/B1 ;
  wire  \picorv32_core/sel38_b1/B2 ;
  wire  \picorv32_core/sel38_b1/B3 ;
  wire  \picorv32_core/sel38_b1/B4 ;
  wire  \picorv32_core/sel38_b1/B5 ;
  wire  \picorv32_core/sel38_b1/B6 ;
  wire  \picorv32_core/sel38_b1/B7 ;
  wire  \picorv32_core/sel38_b2/B0 ;
  wire  \picorv32_core/sel38_b2/B1 ;
  wire  \picorv32_core/sel38_b2/B2 ;
  wire  \picorv32_core/sel38_b2/B3 ;
  wire  \picorv32_core/sel38_b2/B4 ;
  wire  \picorv32_core/sel38_b2/B5 ;
  wire  \picorv32_core/sel38_b2/B6 ;
  wire  \picorv32_core/sel38_b2/B7 ;
  wire  \picorv32_core/sel38_b3/B0 ;
  wire  \picorv32_core/sel38_b3/B1 ;
  wire  \picorv32_core/sel38_b3/B2 ;
  wire  \picorv32_core/sel38_b3/B3 ;
  wire  \picorv32_core/sel38_b3/B4 ;
  wire  \picorv32_core/sel38_b3/B5 ;
  wire  \picorv32_core/sel38_b3/B6 ;
  wire  \picorv32_core/sel38_b3/B7 ;
  wire  \picorv32_core/sel38_b4/B0 ;
  wire  \picorv32_core/sel38_b4/B1 ;
  wire  \picorv32_core/sel38_b4/B2 ;
  wire  \picorv32_core/sel38_b4/B3 ;
  wire  \picorv32_core/sel38_b4/B4 ;
  wire  \picorv32_core/sel38_b4/B5 ;
  wire  \picorv32_core/sel38_b4/B6 ;
  wire  \picorv32_core/sel38_b4/B7 ;
  wire  \picorv32_core/sel40_b0/B0 ;
  wire  \picorv32_core/sel40_b0/B1 ;
  wire  \picorv32_core/sel40_b0/B2 ;
  wire  \picorv32_core/sel40_b0/B3 ;
  wire  \picorv32_core/sel40_b0/B5 ;
  wire  \picorv32_core/sel40_b0/B6 ;
  wire  \picorv32_core/sel40_b0/B7 ;
  wire  \picorv32_core/sel40_b1/B0 ;
  wire  \picorv32_core/sel40_b1/B1 ;
  wire  \picorv32_core/sel40_b1/B2 ;
  wire  \picorv32_core/sel40_b1/B3 ;
  wire  \picorv32_core/sel40_b1/B4 ;
  wire  \picorv32_core/sel40_b1/B5 ;
  wire  \picorv32_core/sel40_b1/B6 ;
  wire  \picorv32_core/sel40_b1/B7 ;
  wire  \picorv32_core/sel40_b2/B0 ;
  wire  \picorv32_core/sel40_b2/B1 ;
  wire  \picorv32_core/sel40_b2/B2 ;
  wire  \picorv32_core/sel40_b2/B3 ;
  wire  \picorv32_core/sel40_b2/B4 ;
  wire  \picorv32_core/sel40_b2/B5 ;
  wire  \picorv32_core/sel40_b2/B6 ;
  wire  \picorv32_core/sel40_b2/B7 ;
  wire  \picorv32_core/sel40_b3/B0 ;
  wire  \picorv32_core/sel40_b3/B1 ;
  wire  \picorv32_core/sel40_b3/B2 ;
  wire  \picorv32_core/sel40_b3/B3 ;
  wire  \picorv32_core/sel40_b3/B4 ;
  wire  \picorv32_core/sel40_b3/B5 ;
  wire  \picorv32_core/sel40_b3/B6 ;
  wire  \picorv32_core/sel40_b3/B7 ;
  wire  \picorv32_core/sel40_b4/B0 ;
  wire  \picorv32_core/sel40_b4/B1 ;
  wire  \picorv32_core/sel40_b4/B2 ;
  wire  \picorv32_core/sel40_b4/B3 ;
  wire  \picorv32_core/sel40_b4/B6 ;
  wire  \picorv32_core/sel40_b4/B7 ;
  wire  \picorv32_core/sel40_b5/B0 ;
  wire  \picorv32_core/sel40_b5/B1 ;
  wire  \picorv32_core/sel40_b5/B2 ;
  wire  \picorv32_core/sel40_b5/B3 ;
  wire  \picorv32_core/sel40_b5/B6 ;
  wire  \picorv32_core/sel40_b5/B7 ;
  wire  \picorv32_core/sel40_b6/B0 ;
  wire  \picorv32_core/sel40_b6/B1 ;
  wire  \picorv32_core/sel40_b6/B2 ;
  wire  \picorv32_core/sel40_b6/B3 ;
  wire  \picorv32_core/sel40_b6/B5 ;
  wire  \picorv32_core/sel40_b6/B6 ;
  wire  \picorv32_core/sel40_b6/B7 ;
  wire  \picorv32_core/sel40_b7/B0 ;
  wire  \picorv32_core/sel40_b7/B1 ;
  wire  \picorv32_core/sel40_b7/B2 ;
  wire  \picorv32_core/sel40_b7/B3 ;
  wire  \picorv32_core/sel40_b7/B5 ;
  wire  \picorv32_core/sel40_b7/B6 ;
  wire  \picorv32_core/sel40_b7/B7 ;
  wire  \picorv32_core/sel41_b0/B0 ;
  wire  \picorv32_core/sel41_b0/B1 ;
  wire  \picorv32_core/sel41_b0/B2 ;
  wire  \picorv32_core/sel41_b0/B3 ;
  wire  \picorv32_core/sel41_b0/B4 ;
  wire  \picorv32_core/sel41_b0/B5 ;
  wire  \picorv32_core/sel41_b0/B6 ;
  wire  \picorv32_core/sel41_b0/B7 ;
  wire  \picorv32_core/sel41_b1/B0 ;
  wire  \picorv32_core/sel41_b1/B1 ;
  wire  \picorv32_core/sel41_b1/B2 ;
  wire  \picorv32_core/sel41_b1/B3 ;
  wire  \picorv32_core/sel41_b1/B4 ;
  wire  \picorv32_core/sel41_b1/B5 ;
  wire  \picorv32_core/sel41_b1/B6 ;
  wire  \picorv32_core/sel41_b1/B7 ;
  wire  \picorv32_core/sel41_b10/B0 ;
  wire  \picorv32_core/sel41_b10/B1 ;
  wire  \picorv32_core/sel41_b10/B2 ;
  wire  \picorv32_core/sel41_b10/B3 ;
  wire  \picorv32_core/sel41_b10/B4 ;
  wire  \picorv32_core/sel41_b10/B5 ;
  wire  \picorv32_core/sel41_b10/B6 ;
  wire  \picorv32_core/sel41_b10/B7 ;
  wire  \picorv32_core/sel41_b11/B0 ;
  wire  \picorv32_core/sel41_b11/B1 ;
  wire  \picorv32_core/sel41_b11/B2 ;
  wire  \picorv32_core/sel41_b11/B3 ;
  wire  \picorv32_core/sel41_b11/B4 ;
  wire  \picorv32_core/sel41_b11/B5 ;
  wire  \picorv32_core/sel41_b11/B6 ;
  wire  \picorv32_core/sel41_b11/B7 ;
  wire  \picorv32_core/sel41_b12/B0 ;
  wire  \picorv32_core/sel41_b12/B1 ;
  wire  \picorv32_core/sel41_b12/B2 ;
  wire  \picorv32_core/sel41_b12/B3 ;
  wire  \picorv32_core/sel41_b12/B4 ;
  wire  \picorv32_core/sel41_b12/B5 ;
  wire  \picorv32_core/sel41_b12/B6 ;
  wire  \picorv32_core/sel41_b12/B7 ;
  wire  \picorv32_core/sel41_b13/B0 ;
  wire  \picorv32_core/sel41_b13/B1 ;
  wire  \picorv32_core/sel41_b13/B2 ;
  wire  \picorv32_core/sel41_b13/B3 ;
  wire  \picorv32_core/sel41_b13/B4 ;
  wire  \picorv32_core/sel41_b13/B5 ;
  wire  \picorv32_core/sel41_b13/B6 ;
  wire  \picorv32_core/sel41_b13/B7 ;
  wire  \picorv32_core/sel41_b14/B0 ;
  wire  \picorv32_core/sel41_b14/B1 ;
  wire  \picorv32_core/sel41_b14/B2 ;
  wire  \picorv32_core/sel41_b14/B3 ;
  wire  \picorv32_core/sel41_b14/B4 ;
  wire  \picorv32_core/sel41_b14/B5 ;
  wire  \picorv32_core/sel41_b14/B6 ;
  wire  \picorv32_core/sel41_b14/B7 ;
  wire  \picorv32_core/sel41_b15/B0 ;
  wire  \picorv32_core/sel41_b15/B1 ;
  wire  \picorv32_core/sel41_b15/B2 ;
  wire  \picorv32_core/sel41_b15/B3 ;
  wire  \picorv32_core/sel41_b15/B4 ;
  wire  \picorv32_core/sel41_b15/B5 ;
  wire  \picorv32_core/sel41_b15/B6 ;
  wire  \picorv32_core/sel41_b15/B7 ;
  wire  \picorv32_core/sel41_b16/B0 ;
  wire  \picorv32_core/sel41_b16/B1 ;
  wire  \picorv32_core/sel41_b16/B2 ;
  wire  \picorv32_core/sel41_b16/B3 ;
  wire  \picorv32_core/sel41_b16/B4 ;
  wire  \picorv32_core/sel41_b16/B5 ;
  wire  \picorv32_core/sel41_b16/B6 ;
  wire  \picorv32_core/sel41_b16/B7 ;
  wire  \picorv32_core/sel41_b17/B0 ;
  wire  \picorv32_core/sel41_b17/B1 ;
  wire  \picorv32_core/sel41_b17/B2 ;
  wire  \picorv32_core/sel41_b17/B3 ;
  wire  \picorv32_core/sel41_b17/B4 ;
  wire  \picorv32_core/sel41_b17/B5 ;
  wire  \picorv32_core/sel41_b17/B6 ;
  wire  \picorv32_core/sel41_b17/B7 ;
  wire  \picorv32_core/sel41_b18/B0 ;
  wire  \picorv32_core/sel41_b18/B1 ;
  wire  \picorv32_core/sel41_b18/B2 ;
  wire  \picorv32_core/sel41_b18/B3 ;
  wire  \picorv32_core/sel41_b18/B4 ;
  wire  \picorv32_core/sel41_b18/B5 ;
  wire  \picorv32_core/sel41_b18/B6 ;
  wire  \picorv32_core/sel41_b18/B7 ;
  wire  \picorv32_core/sel41_b19/B0 ;
  wire  \picorv32_core/sel41_b19/B1 ;
  wire  \picorv32_core/sel41_b19/B2 ;
  wire  \picorv32_core/sel41_b19/B3 ;
  wire  \picorv32_core/sel41_b19/B4 ;
  wire  \picorv32_core/sel41_b19/B5 ;
  wire  \picorv32_core/sel41_b19/B6 ;
  wire  \picorv32_core/sel41_b19/B7 ;
  wire  \picorv32_core/sel41_b2/B0 ;
  wire  \picorv32_core/sel41_b2/B1 ;
  wire  \picorv32_core/sel41_b2/B2 ;
  wire  \picorv32_core/sel41_b2/B3 ;
  wire  \picorv32_core/sel41_b2/B4 ;
  wire  \picorv32_core/sel41_b2/B5 ;
  wire  \picorv32_core/sel41_b2/B6 ;
  wire  \picorv32_core/sel41_b2/B7 ;
  wire  \picorv32_core/sel41_b20/B0 ;
  wire  \picorv32_core/sel41_b20/B1 ;
  wire  \picorv32_core/sel41_b20/B2 ;
  wire  \picorv32_core/sel41_b20/B3 ;
  wire  \picorv32_core/sel41_b20/B4 ;
  wire  \picorv32_core/sel41_b20/B5 ;
  wire  \picorv32_core/sel41_b20/B6 ;
  wire  \picorv32_core/sel41_b20/B7 ;
  wire  \picorv32_core/sel41_b21/B0 ;
  wire  \picorv32_core/sel41_b21/B1 ;
  wire  \picorv32_core/sel41_b21/B2 ;
  wire  \picorv32_core/sel41_b21/B3 ;
  wire  \picorv32_core/sel41_b21/B4 ;
  wire  \picorv32_core/sel41_b21/B5 ;
  wire  \picorv32_core/sel41_b21/B6 ;
  wire  \picorv32_core/sel41_b21/B7 ;
  wire  \picorv32_core/sel41_b22/B0 ;
  wire  \picorv32_core/sel41_b22/B1 ;
  wire  \picorv32_core/sel41_b22/B2 ;
  wire  \picorv32_core/sel41_b22/B3 ;
  wire  \picorv32_core/sel41_b22/B4 ;
  wire  \picorv32_core/sel41_b22/B5 ;
  wire  \picorv32_core/sel41_b22/B6 ;
  wire  \picorv32_core/sel41_b22/B7 ;
  wire  \picorv32_core/sel41_b23/B0 ;
  wire  \picorv32_core/sel41_b23/B1 ;
  wire  \picorv32_core/sel41_b23/B2 ;
  wire  \picorv32_core/sel41_b23/B3 ;
  wire  \picorv32_core/sel41_b23/B4 ;
  wire  \picorv32_core/sel41_b23/B5 ;
  wire  \picorv32_core/sel41_b23/B6 ;
  wire  \picorv32_core/sel41_b23/B7 ;
  wire  \picorv32_core/sel41_b24/B0 ;
  wire  \picorv32_core/sel41_b24/B1 ;
  wire  \picorv32_core/sel41_b24/B2 ;
  wire  \picorv32_core/sel41_b24/B3 ;
  wire  \picorv32_core/sel41_b24/B4 ;
  wire  \picorv32_core/sel41_b24/B5 ;
  wire  \picorv32_core/sel41_b24/B6 ;
  wire  \picorv32_core/sel41_b24/B7 ;
  wire  \picorv32_core/sel41_b25/B0 ;
  wire  \picorv32_core/sel41_b25/B1 ;
  wire  \picorv32_core/sel41_b25/B2 ;
  wire  \picorv32_core/sel41_b25/B3 ;
  wire  \picorv32_core/sel41_b25/B4 ;
  wire  \picorv32_core/sel41_b25/B5 ;
  wire  \picorv32_core/sel41_b25/B6 ;
  wire  \picorv32_core/sel41_b25/B7 ;
  wire  \picorv32_core/sel41_b26/B0 ;
  wire  \picorv32_core/sel41_b26/B1 ;
  wire  \picorv32_core/sel41_b26/B2 ;
  wire  \picorv32_core/sel41_b26/B3 ;
  wire  \picorv32_core/sel41_b26/B4 ;
  wire  \picorv32_core/sel41_b26/B5 ;
  wire  \picorv32_core/sel41_b26/B6 ;
  wire  \picorv32_core/sel41_b26/B7 ;
  wire  \picorv32_core/sel41_b27/B0 ;
  wire  \picorv32_core/sel41_b27/B1 ;
  wire  \picorv32_core/sel41_b27/B2 ;
  wire  \picorv32_core/sel41_b27/B3 ;
  wire  \picorv32_core/sel41_b27/B4 ;
  wire  \picorv32_core/sel41_b27/B5 ;
  wire  \picorv32_core/sel41_b27/B6 ;
  wire  \picorv32_core/sel41_b27/B7 ;
  wire  \picorv32_core/sel41_b28/B0 ;
  wire  \picorv32_core/sel41_b28/B1 ;
  wire  \picorv32_core/sel41_b28/B2 ;
  wire  \picorv32_core/sel41_b28/B3 ;
  wire  \picorv32_core/sel41_b28/B4 ;
  wire  \picorv32_core/sel41_b28/B5 ;
  wire  \picorv32_core/sel41_b28/B6 ;
  wire  \picorv32_core/sel41_b28/B7 ;
  wire  \picorv32_core/sel41_b29/B0 ;
  wire  \picorv32_core/sel41_b29/B1 ;
  wire  \picorv32_core/sel41_b29/B2 ;
  wire  \picorv32_core/sel41_b29/B3 ;
  wire  \picorv32_core/sel41_b29/B4 ;
  wire  \picorv32_core/sel41_b29/B5 ;
  wire  \picorv32_core/sel41_b29/B6 ;
  wire  \picorv32_core/sel41_b29/B7 ;
  wire  \picorv32_core/sel41_b3/B0 ;
  wire  \picorv32_core/sel41_b3/B1 ;
  wire  \picorv32_core/sel41_b3/B2 ;
  wire  \picorv32_core/sel41_b3/B3 ;
  wire  \picorv32_core/sel41_b3/B4 ;
  wire  \picorv32_core/sel41_b3/B5 ;
  wire  \picorv32_core/sel41_b3/B6 ;
  wire  \picorv32_core/sel41_b3/B7 ;
  wire  \picorv32_core/sel41_b30/B0 ;
  wire  \picorv32_core/sel41_b30/B1 ;
  wire  \picorv32_core/sel41_b30/B2 ;
  wire  \picorv32_core/sel41_b30/B3 ;
  wire  \picorv32_core/sel41_b30/B4 ;
  wire  \picorv32_core/sel41_b30/B5 ;
  wire  \picorv32_core/sel41_b30/B6 ;
  wire  \picorv32_core/sel41_b30/B7 ;
  wire  \picorv32_core/sel41_b31/B0 ;
  wire  \picorv32_core/sel41_b31/B1 ;
  wire  \picorv32_core/sel41_b31/B2 ;
  wire  \picorv32_core/sel41_b31/B3 ;
  wire  \picorv32_core/sel41_b31/B4 ;
  wire  \picorv32_core/sel41_b31/B5 ;
  wire  \picorv32_core/sel41_b31/B6 ;
  wire  \picorv32_core/sel41_b31/B7 ;
  wire  \picorv32_core/sel41_b4/B0 ;
  wire  \picorv32_core/sel41_b4/B1 ;
  wire  \picorv32_core/sel41_b4/B2 ;
  wire  \picorv32_core/sel41_b4/B3 ;
  wire  \picorv32_core/sel41_b4/B4 ;
  wire  \picorv32_core/sel41_b4/B5 ;
  wire  \picorv32_core/sel41_b4/B6 ;
  wire  \picorv32_core/sel41_b4/B7 ;
  wire  \picorv32_core/sel41_b5/B0 ;
  wire  \picorv32_core/sel41_b5/B1 ;
  wire  \picorv32_core/sel41_b5/B2 ;
  wire  \picorv32_core/sel41_b5/B3 ;
  wire  \picorv32_core/sel41_b5/B4 ;
  wire  \picorv32_core/sel41_b5/B5 ;
  wire  \picorv32_core/sel41_b5/B6 ;
  wire  \picorv32_core/sel41_b5/B7 ;
  wire  \picorv32_core/sel41_b6/B0 ;
  wire  \picorv32_core/sel41_b6/B1 ;
  wire  \picorv32_core/sel41_b6/B2 ;
  wire  \picorv32_core/sel41_b6/B3 ;
  wire  \picorv32_core/sel41_b6/B4 ;
  wire  \picorv32_core/sel41_b6/B5 ;
  wire  \picorv32_core/sel41_b6/B6 ;
  wire  \picorv32_core/sel41_b6/B7 ;
  wire  \picorv32_core/sel41_b7/B0 ;
  wire  \picorv32_core/sel41_b7/B1 ;
  wire  \picorv32_core/sel41_b7/B2 ;
  wire  \picorv32_core/sel41_b7/B3 ;
  wire  \picorv32_core/sel41_b7/B4 ;
  wire  \picorv32_core/sel41_b7/B5 ;
  wire  \picorv32_core/sel41_b7/B6 ;
  wire  \picorv32_core/sel41_b7/B7 ;
  wire  \picorv32_core/sel41_b8/B0 ;
  wire  \picorv32_core/sel41_b8/B1 ;
  wire  \picorv32_core/sel41_b8/B2 ;
  wire  \picorv32_core/sel41_b8/B3 ;
  wire  \picorv32_core/sel41_b8/B4 ;
  wire  \picorv32_core/sel41_b8/B5 ;
  wire  \picorv32_core/sel41_b8/B6 ;
  wire  \picorv32_core/sel41_b8/B7 ;
  wire  \picorv32_core/sel41_b9/B0 ;
  wire  \picorv32_core/sel41_b9/B1 ;
  wire  \picorv32_core/sel41_b9/B2 ;
  wire  \picorv32_core/sel41_b9/B3 ;
  wire  \picorv32_core/sel41_b9/B4 ;
  wire  \picorv32_core/sel41_b9/B5 ;
  wire  \picorv32_core/sel41_b9/B6 ;
  wire  \picorv32_core/sel41_b9/B7 ;
  wire  \picorv32_core/sel42_b0/B0 ;
  wire  \picorv32_core/sel42_b0/B1 ;
  wire  \picorv32_core/sel42_b0/B2 ;
  wire  \picorv32_core/sel42_b0/B3 ;
  wire  \picorv32_core/sel42_b0/B4 ;
  wire  \picorv32_core/sel42_b0/B5 ;
  wire  \picorv32_core/sel42_b0/B6 ;
  wire  \picorv32_core/sel42_b0/B7 ;
  wire  \picorv32_core/sel42_b1/B0 ;
  wire  \picorv32_core/sel42_b1/B1 ;
  wire  \picorv32_core/sel42_b1/B2 ;
  wire  \picorv32_core/sel42_b1/B3 ;
  wire  \picorv32_core/sel42_b1/B4 ;
  wire  \picorv32_core/sel42_b1/B5 ;
  wire  \picorv32_core/sel42_b1/B6 ;
  wire  \picorv32_core/sel42_b1/B7 ;
  wire  \picorv32_core/sel42_b10/B0 ;
  wire  \picorv32_core/sel42_b10/B1 ;
  wire  \picorv32_core/sel42_b10/B2 ;
  wire  \picorv32_core/sel42_b10/B3 ;
  wire  \picorv32_core/sel42_b10/B4 ;
  wire  \picorv32_core/sel42_b10/B5 ;
  wire  \picorv32_core/sel42_b10/B6 ;
  wire  \picorv32_core/sel42_b10/B7 ;
  wire  \picorv32_core/sel42_b11/B0 ;
  wire  \picorv32_core/sel42_b11/B1 ;
  wire  \picorv32_core/sel42_b11/B2 ;
  wire  \picorv32_core/sel42_b11/B3 ;
  wire  \picorv32_core/sel42_b11/B4 ;
  wire  \picorv32_core/sel42_b11/B5 ;
  wire  \picorv32_core/sel42_b11/B6 ;
  wire  \picorv32_core/sel42_b11/B7 ;
  wire  \picorv32_core/sel42_b12/B0 ;
  wire  \picorv32_core/sel42_b12/B1 ;
  wire  \picorv32_core/sel42_b12/B2 ;
  wire  \picorv32_core/sel42_b12/B3 ;
  wire  \picorv32_core/sel42_b12/B4 ;
  wire  \picorv32_core/sel42_b12/B5 ;
  wire  \picorv32_core/sel42_b12/B6 ;
  wire  \picorv32_core/sel42_b12/B7 ;
  wire  \picorv32_core/sel42_b13/B0 ;
  wire  \picorv32_core/sel42_b13/B1 ;
  wire  \picorv32_core/sel42_b13/B2 ;
  wire  \picorv32_core/sel42_b13/B3 ;
  wire  \picorv32_core/sel42_b13/B4 ;
  wire  \picorv32_core/sel42_b13/B5 ;
  wire  \picorv32_core/sel42_b13/B6 ;
  wire  \picorv32_core/sel42_b13/B7 ;
  wire  \picorv32_core/sel42_b14/B0 ;
  wire  \picorv32_core/sel42_b14/B1 ;
  wire  \picorv32_core/sel42_b14/B2 ;
  wire  \picorv32_core/sel42_b14/B3 ;
  wire  \picorv32_core/sel42_b14/B4 ;
  wire  \picorv32_core/sel42_b14/B5 ;
  wire  \picorv32_core/sel42_b14/B6 ;
  wire  \picorv32_core/sel42_b14/B7 ;
  wire  \picorv32_core/sel42_b15/B0 ;
  wire  \picorv32_core/sel42_b15/B1 ;
  wire  \picorv32_core/sel42_b15/B2 ;
  wire  \picorv32_core/sel42_b15/B3 ;
  wire  \picorv32_core/sel42_b15/B4 ;
  wire  \picorv32_core/sel42_b15/B5 ;
  wire  \picorv32_core/sel42_b15/B6 ;
  wire  \picorv32_core/sel42_b15/B7 ;
  wire  \picorv32_core/sel42_b16/B0 ;
  wire  \picorv32_core/sel42_b16/B1 ;
  wire  \picorv32_core/sel42_b16/B2 ;
  wire  \picorv32_core/sel42_b16/B3 ;
  wire  \picorv32_core/sel42_b16/B4 ;
  wire  \picorv32_core/sel42_b16/B5 ;
  wire  \picorv32_core/sel42_b16/B6 ;
  wire  \picorv32_core/sel42_b16/B7 ;
  wire  \picorv32_core/sel42_b17/B0 ;
  wire  \picorv32_core/sel42_b17/B1 ;
  wire  \picorv32_core/sel42_b17/B2 ;
  wire  \picorv32_core/sel42_b17/B3 ;
  wire  \picorv32_core/sel42_b17/B4 ;
  wire  \picorv32_core/sel42_b17/B5 ;
  wire  \picorv32_core/sel42_b17/B6 ;
  wire  \picorv32_core/sel42_b17/B7 ;
  wire  \picorv32_core/sel42_b18/B0 ;
  wire  \picorv32_core/sel42_b18/B1 ;
  wire  \picorv32_core/sel42_b18/B2 ;
  wire  \picorv32_core/sel42_b18/B3 ;
  wire  \picorv32_core/sel42_b18/B4 ;
  wire  \picorv32_core/sel42_b18/B5 ;
  wire  \picorv32_core/sel42_b18/B6 ;
  wire  \picorv32_core/sel42_b18/B7 ;
  wire  \picorv32_core/sel42_b19/B0 ;
  wire  \picorv32_core/sel42_b19/B1 ;
  wire  \picorv32_core/sel42_b19/B2 ;
  wire  \picorv32_core/sel42_b19/B3 ;
  wire  \picorv32_core/sel42_b19/B4 ;
  wire  \picorv32_core/sel42_b19/B5 ;
  wire  \picorv32_core/sel42_b19/B6 ;
  wire  \picorv32_core/sel42_b19/B7 ;
  wire  \picorv32_core/sel42_b2/B0 ;
  wire  \picorv32_core/sel42_b2/B1 ;
  wire  \picorv32_core/sel42_b2/B2 ;
  wire  \picorv32_core/sel42_b2/B3 ;
  wire  \picorv32_core/sel42_b2/B4 ;
  wire  \picorv32_core/sel42_b2/B5 ;
  wire  \picorv32_core/sel42_b2/B6 ;
  wire  \picorv32_core/sel42_b2/B7 ;
  wire  \picorv32_core/sel42_b20/B0 ;
  wire  \picorv32_core/sel42_b20/B1 ;
  wire  \picorv32_core/sel42_b20/B2 ;
  wire  \picorv32_core/sel42_b20/B3 ;
  wire  \picorv32_core/sel42_b20/B4 ;
  wire  \picorv32_core/sel42_b20/B5 ;
  wire  \picorv32_core/sel42_b20/B6 ;
  wire  \picorv32_core/sel42_b20/B7 ;
  wire  \picorv32_core/sel42_b21/B0 ;
  wire  \picorv32_core/sel42_b21/B1 ;
  wire  \picorv32_core/sel42_b21/B2 ;
  wire  \picorv32_core/sel42_b21/B3 ;
  wire  \picorv32_core/sel42_b21/B4 ;
  wire  \picorv32_core/sel42_b21/B5 ;
  wire  \picorv32_core/sel42_b21/B6 ;
  wire  \picorv32_core/sel42_b21/B7 ;
  wire  \picorv32_core/sel42_b22/B0 ;
  wire  \picorv32_core/sel42_b22/B1 ;
  wire  \picorv32_core/sel42_b22/B2 ;
  wire  \picorv32_core/sel42_b22/B3 ;
  wire  \picorv32_core/sel42_b22/B4 ;
  wire  \picorv32_core/sel42_b22/B5 ;
  wire  \picorv32_core/sel42_b22/B6 ;
  wire  \picorv32_core/sel42_b22/B7 ;
  wire  \picorv32_core/sel42_b23/B0 ;
  wire  \picorv32_core/sel42_b23/B1 ;
  wire  \picorv32_core/sel42_b23/B2 ;
  wire  \picorv32_core/sel42_b23/B3 ;
  wire  \picorv32_core/sel42_b23/B4 ;
  wire  \picorv32_core/sel42_b23/B5 ;
  wire  \picorv32_core/sel42_b23/B6 ;
  wire  \picorv32_core/sel42_b23/B7 ;
  wire  \picorv32_core/sel42_b24/B0 ;
  wire  \picorv32_core/sel42_b24/B1 ;
  wire  \picorv32_core/sel42_b24/B2 ;
  wire  \picorv32_core/sel42_b24/B3 ;
  wire  \picorv32_core/sel42_b24/B4 ;
  wire  \picorv32_core/sel42_b24/B5 ;
  wire  \picorv32_core/sel42_b24/B6 ;
  wire  \picorv32_core/sel42_b24/B7 ;
  wire  \picorv32_core/sel42_b25/B0 ;
  wire  \picorv32_core/sel42_b25/B1 ;
  wire  \picorv32_core/sel42_b25/B2 ;
  wire  \picorv32_core/sel42_b25/B3 ;
  wire  \picorv32_core/sel42_b25/B4 ;
  wire  \picorv32_core/sel42_b25/B5 ;
  wire  \picorv32_core/sel42_b25/B6 ;
  wire  \picorv32_core/sel42_b25/B7 ;
  wire  \picorv32_core/sel42_b26/B0 ;
  wire  \picorv32_core/sel42_b26/B1 ;
  wire  \picorv32_core/sel42_b26/B2 ;
  wire  \picorv32_core/sel42_b26/B3 ;
  wire  \picorv32_core/sel42_b26/B4 ;
  wire  \picorv32_core/sel42_b26/B5 ;
  wire  \picorv32_core/sel42_b26/B6 ;
  wire  \picorv32_core/sel42_b26/B7 ;
  wire  \picorv32_core/sel42_b27/B0 ;
  wire  \picorv32_core/sel42_b27/B1 ;
  wire  \picorv32_core/sel42_b27/B2 ;
  wire  \picorv32_core/sel42_b27/B3 ;
  wire  \picorv32_core/sel42_b27/B4 ;
  wire  \picorv32_core/sel42_b27/B5 ;
  wire  \picorv32_core/sel42_b27/B6 ;
  wire  \picorv32_core/sel42_b27/B7 ;
  wire  \picorv32_core/sel42_b28/B0 ;
  wire  \picorv32_core/sel42_b28/B1 ;
  wire  \picorv32_core/sel42_b28/B2 ;
  wire  \picorv32_core/sel42_b28/B3 ;
  wire  \picorv32_core/sel42_b28/B4 ;
  wire  \picorv32_core/sel42_b28/B5 ;
  wire  \picorv32_core/sel42_b28/B6 ;
  wire  \picorv32_core/sel42_b28/B7 ;
  wire  \picorv32_core/sel42_b29/B0 ;
  wire  \picorv32_core/sel42_b29/B1 ;
  wire  \picorv32_core/sel42_b29/B2 ;
  wire  \picorv32_core/sel42_b29/B3 ;
  wire  \picorv32_core/sel42_b29/B4 ;
  wire  \picorv32_core/sel42_b29/B5 ;
  wire  \picorv32_core/sel42_b29/B6 ;
  wire  \picorv32_core/sel42_b29/B7 ;
  wire  \picorv32_core/sel42_b3/B0 ;
  wire  \picorv32_core/sel42_b3/B1 ;
  wire  \picorv32_core/sel42_b3/B2 ;
  wire  \picorv32_core/sel42_b3/B3 ;
  wire  \picorv32_core/sel42_b3/B4 ;
  wire  \picorv32_core/sel42_b3/B5 ;
  wire  \picorv32_core/sel42_b3/B6 ;
  wire  \picorv32_core/sel42_b3/B7 ;
  wire  \picorv32_core/sel42_b30/B0 ;
  wire  \picorv32_core/sel42_b30/B1 ;
  wire  \picorv32_core/sel42_b30/B2 ;
  wire  \picorv32_core/sel42_b30/B3 ;
  wire  \picorv32_core/sel42_b30/B4 ;
  wire  \picorv32_core/sel42_b30/B5 ;
  wire  \picorv32_core/sel42_b30/B6 ;
  wire  \picorv32_core/sel42_b30/B7 ;
  wire  \picorv32_core/sel42_b31/B0 ;
  wire  \picorv32_core/sel42_b31/B1 ;
  wire  \picorv32_core/sel42_b31/B2 ;
  wire  \picorv32_core/sel42_b31/B3 ;
  wire  \picorv32_core/sel42_b31/B4 ;
  wire  \picorv32_core/sel42_b31/B5 ;
  wire  \picorv32_core/sel42_b31/B6 ;
  wire  \picorv32_core/sel42_b31/B7 ;
  wire  \picorv32_core/sel42_b4/B0 ;
  wire  \picorv32_core/sel42_b4/B1 ;
  wire  \picorv32_core/sel42_b4/B2 ;
  wire  \picorv32_core/sel42_b4/B3 ;
  wire  \picorv32_core/sel42_b4/B4 ;
  wire  \picorv32_core/sel42_b4/B5 ;
  wire  \picorv32_core/sel42_b4/B6 ;
  wire  \picorv32_core/sel42_b4/B7 ;
  wire  \picorv32_core/sel42_b5/B0 ;
  wire  \picorv32_core/sel42_b5/B1 ;
  wire  \picorv32_core/sel42_b5/B2 ;
  wire  \picorv32_core/sel42_b5/B3 ;
  wire  \picorv32_core/sel42_b5/B4 ;
  wire  \picorv32_core/sel42_b5/B5 ;
  wire  \picorv32_core/sel42_b5/B6 ;
  wire  \picorv32_core/sel42_b5/B7 ;
  wire  \picorv32_core/sel42_b6/B0 ;
  wire  \picorv32_core/sel42_b6/B1 ;
  wire  \picorv32_core/sel42_b6/B2 ;
  wire  \picorv32_core/sel42_b6/B3 ;
  wire  \picorv32_core/sel42_b6/B4 ;
  wire  \picorv32_core/sel42_b6/B5 ;
  wire  \picorv32_core/sel42_b6/B6 ;
  wire  \picorv32_core/sel42_b6/B7 ;
  wire  \picorv32_core/sel42_b7/B0 ;
  wire  \picorv32_core/sel42_b7/B1 ;
  wire  \picorv32_core/sel42_b7/B2 ;
  wire  \picorv32_core/sel42_b7/B3 ;
  wire  \picorv32_core/sel42_b7/B4 ;
  wire  \picorv32_core/sel42_b7/B5 ;
  wire  \picorv32_core/sel42_b7/B6 ;
  wire  \picorv32_core/sel42_b7/B7 ;
  wire  \picorv32_core/sel42_b8/B0 ;
  wire  \picorv32_core/sel42_b8/B1 ;
  wire  \picorv32_core/sel42_b8/B2 ;
  wire  \picorv32_core/sel42_b8/B3 ;
  wire  \picorv32_core/sel42_b8/B4 ;
  wire  \picorv32_core/sel42_b8/B5 ;
  wire  \picorv32_core/sel42_b8/B6 ;
  wire  \picorv32_core/sel42_b8/B7 ;
  wire  \picorv32_core/sel42_b9/B0 ;
  wire  \picorv32_core/sel42_b9/B1 ;
  wire  \picorv32_core/sel42_b9/B2 ;
  wire  \picorv32_core/sel42_b9/B3 ;
  wire  \picorv32_core/sel42_b9/B4 ;
  wire  \picorv32_core/sel42_b9/B5 ;
  wire  \picorv32_core/sel42_b9/B6 ;
  wire  \picorv32_core/sel42_b9/B7 ;
  wire  \picorv32_core/sel43_b0/B0 ;
  wire  \picorv32_core/sel43_b0/B2 ;
  wire  \picorv32_core/sel43_b0/B3 ;
  wire  \picorv32_core/sel43_b0/B5 ;
  wire  \picorv32_core/sel43_b1/B0 ;
  wire  \picorv32_core/sel43_b1/B2 ;
  wire  \picorv32_core/sel43_b1/B3 ;
  wire  \picorv32_core/sel43_b1/B5 ;
  wire  \picorv32_core/sel43_b10/B0 ;
  wire  \picorv32_core/sel43_b10/B2 ;
  wire  \picorv32_core/sel43_b10/B3 ;
  wire  \picorv32_core/sel43_b10/B5 ;
  wire  \picorv32_core/sel43_b11/B0 ;
  wire  \picorv32_core/sel43_b11/B2 ;
  wire  \picorv32_core/sel43_b11/B3 ;
  wire  \picorv32_core/sel43_b11/B5 ;
  wire  \picorv32_core/sel43_b12/B0 ;
  wire  \picorv32_core/sel43_b12/B2 ;
  wire  \picorv32_core/sel43_b12/B3 ;
  wire  \picorv32_core/sel43_b12/B5 ;
  wire  \picorv32_core/sel43_b13/B0 ;
  wire  \picorv32_core/sel43_b13/B2 ;
  wire  \picorv32_core/sel43_b13/B3 ;
  wire  \picorv32_core/sel43_b13/B5 ;
  wire  \picorv32_core/sel43_b14/B0 ;
  wire  \picorv32_core/sel43_b14/B2 ;
  wire  \picorv32_core/sel43_b14/B3 ;
  wire  \picorv32_core/sel43_b14/B5 ;
  wire  \picorv32_core/sel43_b15/B0 ;
  wire  \picorv32_core/sel43_b15/B2 ;
  wire  \picorv32_core/sel43_b15/B3 ;
  wire  \picorv32_core/sel43_b15/B5 ;
  wire  \picorv32_core/sel43_b16/B0 ;
  wire  \picorv32_core/sel43_b16/B2 ;
  wire  \picorv32_core/sel43_b16/B3 ;
  wire  \picorv32_core/sel43_b16/B5 ;
  wire  \picorv32_core/sel43_b17/B0 ;
  wire  \picorv32_core/sel43_b17/B2 ;
  wire  \picorv32_core/sel43_b17/B3 ;
  wire  \picorv32_core/sel43_b17/B5 ;
  wire  \picorv32_core/sel43_b18/B0 ;
  wire  \picorv32_core/sel43_b18/B2 ;
  wire  \picorv32_core/sel43_b18/B3 ;
  wire  \picorv32_core/sel43_b18/B5 ;
  wire  \picorv32_core/sel43_b19/B0 ;
  wire  \picorv32_core/sel43_b19/B2 ;
  wire  \picorv32_core/sel43_b19/B3 ;
  wire  \picorv32_core/sel43_b19/B5 ;
  wire  \picorv32_core/sel43_b2/B0 ;
  wire  \picorv32_core/sel43_b2/B2 ;
  wire  \picorv32_core/sel43_b2/B3 ;
  wire  \picorv32_core/sel43_b2/B5 ;
  wire  \picorv32_core/sel43_b20/B0 ;
  wire  \picorv32_core/sel43_b20/B2 ;
  wire  \picorv32_core/sel43_b20/B3 ;
  wire  \picorv32_core/sel43_b20/B5 ;
  wire  \picorv32_core/sel43_b21/B0 ;
  wire  \picorv32_core/sel43_b21/B2 ;
  wire  \picorv32_core/sel43_b21/B3 ;
  wire  \picorv32_core/sel43_b21/B5 ;
  wire  \picorv32_core/sel43_b22/B0 ;
  wire  \picorv32_core/sel43_b22/B2 ;
  wire  \picorv32_core/sel43_b22/B3 ;
  wire  \picorv32_core/sel43_b22/B5 ;
  wire  \picorv32_core/sel43_b23/B0 ;
  wire  \picorv32_core/sel43_b23/B2 ;
  wire  \picorv32_core/sel43_b23/B3 ;
  wire  \picorv32_core/sel43_b23/B5 ;
  wire  \picorv32_core/sel43_b24/B0 ;
  wire  \picorv32_core/sel43_b24/B2 ;
  wire  \picorv32_core/sel43_b24/B3 ;
  wire  \picorv32_core/sel43_b24/B5 ;
  wire  \picorv32_core/sel43_b25/B0 ;
  wire  \picorv32_core/sel43_b25/B2 ;
  wire  \picorv32_core/sel43_b25/B3 ;
  wire  \picorv32_core/sel43_b25/B5 ;
  wire  \picorv32_core/sel43_b26/B0 ;
  wire  \picorv32_core/sel43_b26/B2 ;
  wire  \picorv32_core/sel43_b26/B3 ;
  wire  \picorv32_core/sel43_b26/B5 ;
  wire  \picorv32_core/sel43_b27/B0 ;
  wire  \picorv32_core/sel43_b27/B2 ;
  wire  \picorv32_core/sel43_b27/B3 ;
  wire  \picorv32_core/sel43_b27/B5 ;
  wire  \picorv32_core/sel43_b28/B0 ;
  wire  \picorv32_core/sel43_b28/B2 ;
  wire  \picorv32_core/sel43_b28/B3 ;
  wire  \picorv32_core/sel43_b28/B5 ;
  wire  \picorv32_core/sel43_b29/B0 ;
  wire  \picorv32_core/sel43_b29/B2 ;
  wire  \picorv32_core/sel43_b29/B3 ;
  wire  \picorv32_core/sel43_b29/B5 ;
  wire  \picorv32_core/sel43_b3/B0 ;
  wire  \picorv32_core/sel43_b3/B2 ;
  wire  \picorv32_core/sel43_b3/B3 ;
  wire  \picorv32_core/sel43_b3/B5 ;
  wire  \picorv32_core/sel43_b30/B0 ;
  wire  \picorv32_core/sel43_b30/B2 ;
  wire  \picorv32_core/sel43_b30/B3 ;
  wire  \picorv32_core/sel43_b30/B5 ;
  wire  \picorv32_core/sel43_b31/B0 ;
  wire  \picorv32_core/sel43_b31/B2 ;
  wire  \picorv32_core/sel43_b31/B3 ;
  wire  \picorv32_core/sel43_b31/B5 ;
  wire  \picorv32_core/sel43_b4/B0 ;
  wire  \picorv32_core/sel43_b4/B2 ;
  wire  \picorv32_core/sel43_b4/B3 ;
  wire  \picorv32_core/sel43_b4/B5 ;
  wire  \picorv32_core/sel43_b5/B0 ;
  wire  \picorv32_core/sel43_b5/B2 ;
  wire  \picorv32_core/sel43_b5/B3 ;
  wire  \picorv32_core/sel43_b5/B5 ;
  wire  \picorv32_core/sel43_b6/B0 ;
  wire  \picorv32_core/sel43_b6/B2 ;
  wire  \picorv32_core/sel43_b6/B3 ;
  wire  \picorv32_core/sel43_b6/B5 ;
  wire  \picorv32_core/sel43_b7/B0 ;
  wire  \picorv32_core/sel43_b7/B2 ;
  wire  \picorv32_core/sel43_b7/B3 ;
  wire  \picorv32_core/sel43_b7/B5 ;
  wire  \picorv32_core/sel43_b8/B0 ;
  wire  \picorv32_core/sel43_b8/B2 ;
  wire  \picorv32_core/sel43_b8/B3 ;
  wire  \picorv32_core/sel43_b8/B5 ;
  wire  \picorv32_core/sel43_b9/B0 ;
  wire  \picorv32_core/sel43_b9/B2 ;
  wire  \picorv32_core/sel43_b9/B3 ;
  wire  \picorv32_core/sel43_b9/B5 ;
  wire  \picorv32_core/sel44_b0/B2 ;
  wire  \picorv32_core/sel44_b0/B5 ;
  wire  \picorv32_core/sel44_b1/B2 ;
  wire  \picorv32_core/sel44_b1/B5 ;
  wire  \picorv32_core/sel44_b2/B2 ;
  wire  \picorv32_core/sel44_b2/B5 ;
  wire  \picorv32_core/sel44_b3/B2 ;
  wire  \picorv32_core/sel44_b3/B5 ;
  wire  \picorv32_core/sel44_b4/B2 ;
  wire  \picorv32_core/sel44_b4/B5 ;
  wire  \picorv32_core/sel45/B0 ;
  wire  \picorv32_core/sel45/B1 ;
  wire  \picorv32_core/sel45/B2 ;
  wire  \picorv32_core/sel45/B3 ;
  wire  \picorv32_core/sel4_b0/B0 ;
  wire  \picorv32_core/sel4_b0/B1 ;
  wire  \picorv32_core/sel4_b1/B0 ;
  wire  \picorv32_core/sel4_b1/B1 ;
  wire  \picorv32_core/sel4_b2/B0 ;
  wire  \picorv32_core/sel4_b2/B1 ;
  wire  \picorv32_core/sel4_b2/B2 ;
  wire  \picorv32_core/sel5_b0/B0 ;
  wire  \picorv32_core/sel5_b0/B2 ;
  wire  \picorv32_core/sel5_b1/B0 ;
  wire  \picorv32_core/sel5_b1/B2 ;
  wire  \picorv32_core/sel5_b2/B0 ;
  wire  \picorv32_core/sel5_b2/B1 ;
  wire  \picorv32_core/sel5_b2/B2 ;
  wire  \picorv32_core/sel5_b3/B0 ;
  wire  \picorv32_core/sel5_b3/B1 ;
  wire  \picorv32_core/sel5_b3/B2 ;
  wire  \picorv32_core/sel5_b4/B0 ;
  wire  \picorv32_core/sel5_b4/B1 ;
  wire  \picorv32_core/sel5_b4/B2 ;
  wire  \picorv32_core/sel6_b0/B0 ;
  wire  \picorv32_core/sel6_b1/B0 ;
  wire  \picorv32_core/sel6_b1/B1 ;
  wire  \picorv32_core/sel6_b1/B2 ;
  wire  \picorv32_core/sel6_b2/B0 ;
  wire  \picorv32_core/sel6_b2/B2 ;
  wire  \picorv32_core/sel6_b3/B0 ;
  wire  \picorv32_core/sel6_b3/B2 ;
  wire  \picorv32_core/sel6_b4/B0 ;
  wire  \picorv32_core/sel6_b4/B2 ;
  wire  \picorv32_core/sel7/B1 ;
  wire [3:0] \uart/n100 ;
  wire [3:0] \uart/n101 ;
  wire [2:0] \uart/n102 ;
  wire [7:0] \uart/n106 ;
  wire [31:0] \uart/n16 ;
  wire [3:0] \uart/n31 ;
  wire [3:0] \uart/n32 ;
  wire [4:0] \uart/n33 ;
  wire [3:0] \uart/n35 ;
  wire [3:0] \uart/n36 ;
  wire [3:0] \uart/n37 ;
  wire [3:0] \uart/n38 ;
  wire [3:0] \uart/n4 ;
  wire [7:0] \uart/n45 ;
  wire [2:0] \uart/n46 ;
  wire [3:0] \uart/n47 ;
  wire [3:0] \uart/n48 ;
  wire [3:0] \uart/n49 ;
  wire [31:0] \uart/n5 ;
  wire [3:0] \uart/n50 ;
  wire [3:0] \uart/n54 ;
  wire [3:0] \uart/n55 ;
  wire [4:0] \uart/n57 ;
  wire [7:0] \uart/n59 ;
  wire [31:0] \uart/n6 ;
  wire [1:0] \uart/n61 ;
  wire [1:0] \uart/n63 ;
  wire [1:0] \uart/n65 ;
  wire [1:0] \uart/n67 ;
  wire [1:0] \uart/n69 ;
  wire [1:0] \uart/n71 ;
  wire [1:0] \uart/n73 ;
  wire [1:0] \uart/n75 ;
  wire [7:0] \uart/n76 ;
  wire [3:0] \uart/n77 ;
  wire [7:0] \uart/n78 ;
  wire [3:0] \uart/n79 ;
  wire [3:0] \uart/n80 ;
  wire [3:0] \uart/n81 ;
  wire [3:0] \uart/n92 ;
  wire [31:0] \uart/uart_bsrr ;  // ../src/uart.v(28)
  wire [2:0] \uart/uart_cnt_rx ;  // ../src/uart.v(151)
  wire [31:0] \uart/uart_counter ;  // ../src/uart.v(30)
  wire [7:0] \uart/uart_idr ;  // ../src/uart.v(27)
  wire [7:0] \uart/uart_idr_t ;  // ../src/uart.v(153)
  wire [7:0] \uart/uart_odr ;  // ../src/uart.v(26)
  wire [2:0] \uart/uart_op_clock_by_3_c ;  // ../src/uart.v(35)
  wire [3:0] \uart/uart_smp_rx ;  // ../src/uart.v(152)
  wire [7:0] \uart/uart_sr ;  // ../src/uart.v(42)
  wire [3:0] \uart/uart_status_rxd ;  // ../src/uart.v(148)
  wire [3:0] \uart/uart_status_txd ;  // ../src/uart.v(32)
  wire [31:0] uart_do;  // ../src/top.v(98)
  wire mem_la_addr$2$_neg;
  wire mem_la_addr$3$_neg;
  wire mem_la_write;  // ../src/top.v(28)
  wire mem_la_write_neg;
  wire n0;
  wire n1;
  wire n11;
  wire n13;
  wire n15;
  wire n16;
  wire n2;
  wire n6;
  wire n7;
  wire n9;
  wire \picorv32_core/alu_eq ;  // ../src/picorv32.v(1180)
  wire \picorv32_core/alu_lts ;  // ../src/picorv32.v(1180)
  wire \picorv32_core/alu_ltu ;  // ../src/picorv32.v(1180)
  wire \picorv32_core/alu_out_0 ;  // ../src/picorv32.v(1175)
  wire \picorv32_core/clear_prefetched_high_word ;  // ../src/picorv32.v(330)
  wire \picorv32_core/clear_prefetched_high_word_neg ;
  wire \picorv32_core/clear_prefetched_high_word_q ;  // ../src/picorv32.v(1240)
  wire \picorv32_core/compressed_instr ;  // ../src/picorv32.v(625)
  wire \picorv32_core/cpuregs_write ;  // ../src/picorv32.v(1251)
  wire \picorv32_core/decoder_pseudo_trigger ;  // ../src/picorv32.v(623)
  wire \picorv32_core/decoder_trigger ;  // ../src/picorv32.v(621)
  wire \picorv32_core/instr_add ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_addi ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_and ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_andi ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_auipc ;  // ../src/picorv32.v(610)
  wire \picorv32_core/instr_beq ;  // ../src/picorv32.v(611)
  wire \picorv32_core/instr_bge ;  // ../src/picorv32.v(611)
  wire \picorv32_core/instr_bgeu ;  // ../src/picorv32.v(611)
  wire \picorv32_core/instr_blt ;  // ../src/picorv32.v(611)
  wire \picorv32_core/instr_bltu ;  // ../src/picorv32.v(611)
  wire \picorv32_core/instr_bne ;  // ../src/picorv32.v(611)
  wire \picorv32_core/instr_jal ;  // ../src/picorv32.v(610)
  wire \picorv32_core/instr_jal_neg ;
  wire \picorv32_core/instr_jalr ;  // ../src/picorv32.v(610)
  wire \picorv32_core/instr_lb ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_lbu ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_lh ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_lhu ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_lui ;  // ../src/picorv32.v(610)
  wire \picorv32_core/instr_lw ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_or ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_ori ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_rdcycle ;  // ../src/picorv32.v(615)
  wire \picorv32_core/instr_rdcycleh ;  // ../src/picorv32.v(615)
  wire \picorv32_core/instr_rdinstr ;  // ../src/picorv32.v(615)
  wire \picorv32_core/instr_rdinstrh ;  // ../src/picorv32.v(615)
  wire \picorv32_core/instr_sb ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_sh ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_sll ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_slli ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_slt ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_slti ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_sltiu ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_sltu ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_sra ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_srai ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_srl ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_srli ;  // ../src/picorv32.v(613)
  wire \picorv32_core/instr_sub ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_sw ;  // ../src/picorv32.v(612)
  wire \picorv32_core/instr_trap ;  // ../src/picorv32.v(617)
  wire \picorv32_core/instr_xor ;  // ../src/picorv32.v(614)
  wire \picorv32_core/instr_xori ;  // ../src/picorv32.v(613)
  wire \picorv32_core/is_alu_reg_imm ;  // ../src/picorv32.v(638)
  wire \picorv32_core/is_alu_reg_reg ;  // ../src/picorv32.v(639)
  wire \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ;  // ../src/picorv32.v(636)
  wire \picorv32_core/is_compare ;  // ../src/picorv32.v(640)
  wire \picorv32_core/is_jalr_addi_slti_sltiu_xori_ori_andi ;  // ../src/picorv32.v(630)
  wire \picorv32_core/is_lb_lh_lw_lbu_lhu ;  // ../src/picorv32.v(628)
  wire \picorv32_core/is_lbu_lhu_lw ;  // ../src/picorv32.v(637)
  wire \picorv32_core/is_lui_auipc_jal ;  // ../src/picorv32.v(627)
  wire \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub ;  // ../src/picorv32.v(633)
  wire \picorv32_core/is_rdcycle_rdcycleh_rdinstr_rdinstrh ;  // ../src/picorv32.v(650)
  wire \picorv32_core/is_sb_sh_sw ;  // ../src/picorv32.v(631)
  wire \picorv32_core/is_sll_srl_sra ;  // ../src/picorv32.v(632)
  wire \picorv32_core/is_slli_srli_srai ;  // ../src/picorv32.v(629)
  wire \picorv32_core/is_slti_blt_slt ;  // ../src/picorv32.v(634)
  wire \picorv32_core/is_sltiu_bltu_sltu ;  // ../src/picorv32.v(635)
  wire \picorv32_core/latched_branch ;  // ../src/picorv32.v(1157)
  wire \picorv32_core/latched_compr ;  // ../src/picorv32.v(1158)
  wire \picorv32_core/latched_is_lb ;  // ../src/picorv32.v(1162)
  wire \picorv32_core/latched_is_lh ;  // ../src/picorv32.v(1161)
  wire \picorv32_core/latched_is_lu ;  // ../src/picorv32.v(1160)
  wire \picorv32_core/latched_stalu ;  // ../src/picorv32.v(1156)
  wire \picorv32_core/latched_store ;  // ../src/picorv32.v(1155)
  wire \picorv32_core/mem_do_prefetch ;  // ../src/picorv32.v(320)
  wire \picorv32_core/mem_do_rdata ;  // ../src/picorv32.v(322)
  wire \picorv32_core/mem_do_rinst ;  // ../src/picorv32.v(321)
  wire \picorv32_core/mem_do_wdata ;  // ../src/picorv32.v(323)
  wire \picorv32_core/mem_done ;  // ../src/picorv32.v(340)
  wire \picorv32_core/mem_done_neg ;
  wire \picorv32_core/mem_la_firstword ;  // ../src/picorv32.v(326)
  wire \picorv32_core/mem_la_firstword_neg ;
  wire \picorv32_core/mem_la_firstword_xfer ;  // ../src/picorv32.v(327)
  wire \picorv32_core/mem_la_read ;  // ../src/picorv32.v(87)
  wire \picorv32_core/mem_la_read_neg ;
  wire \picorv32_core/mem_la_secondword ;  // ../src/picorv32.v(325)
  wire \picorv32_core/mem_la_secondword_neg ;
  wire \picorv32_core/mem_la_use_prefetched_high_word ;  // ../src/picorv32.v(336)
  wire \picorv32_core/mem_la_use_prefetched_high_word_neg ;
  wire \picorv32_core/mem_rdata_latched$0$_neg ;
  wire \picorv32_core/mem_rdata_latched$1$_neg ;
  wire \picorv32_core/mem_rdata_latched$13$_neg ;
  wire \picorv32_core/mem_rdata_latched$14$_neg ;
  wire \picorv32_core/mem_rdata_latched$15$_neg ;
  wire \picorv32_core/mem_state$1$_neg ;
  wire \picorv32_core/mem_valid ;  // ../src/picorv32.v(77)
  wire \picorv32_core/mem_wordsize$0$_neg ;
  wire \picorv32_core/mem_wordsize$1$_neg ;
  wire \picorv32_core/mem_xfer ;  // ../src/picorv32.v(337)
  wire \picorv32_core/mux100_sel_is_6_o ;
  wire \picorv32_core/mux103_sel_is_5_o ;
  wire \picorv32_core/mux104_sel_is_5_o ;
  wire \picorv32_core/mux105_sel_is_5_o ;
  wire \picorv32_core/mux127_b0_sel_is_1_o ;
  wire \picorv32_core/mux12_b0_sel_is_3_o ;
  wire \picorv32_core/mux131_b0_sel_is_1_o ;
  wire \picorv32_core/mux132_b0_sel_is_3_o ;
  wire \picorv32_core/mux132_b32_sel_is_3_o ;
  wire \picorv32_core/mux13_b1_sel_is_0_o ;
  wire \picorv32_core/mux13_b2_sel_is_2_o ;
  wire \picorv32_core/mux148_b0_sel_is_3_o ;
  wire \picorv32_core/mux15_b0_sel_is_0_o ;
  wire \picorv32_core/mux162_b0_sel_is_0_o ;
  wire \picorv32_core/mux162_b0_sel_is_0_o_neg ;
  wire \picorv32_core/mux163_b0_sel_is_1_o ;
  wire \picorv32_core/mux163_b0_sel_is_1_o_neg ;
  wire \picorv32_core/mux164_b0_sel_is_0_o ;
  wire \picorv32_core/mux165_b0_sel_is_0_o ;
  wire \picorv32_core/mux19_b0_sel_is_0_o ;
  wire \picorv32_core/mux20_b0_sel_is_2_o ;
  wire \picorv32_core/mux20_b2_sel_is_0_o ;
  wire \picorv32_core/mux21_b0_sel_is_2_o ;
  wire \picorv32_core/mux24_b3_sel_is_3_o ;
  wire \picorv32_core/mux28_b0_sel_is_0_o ;
  wire \picorv32_core/mux32_b0_sel_is_2_o ;
  wire \picorv32_core/mux35_b0_sel_is_2_o ;
  wire \picorv32_core/mux38_b0_sel_is_0_o ;
  wire \picorv32_core/mux3_b16_sel_is_0_o ;
  wire \picorv32_core/mux4_b0_sel_is_0_o ;
  wire \picorv32_core/mux51_b0_sel_is_3_o ;
  wire \picorv32_core/mux55_b10_sel_is_3_o ;
  wire \picorv32_core/mux59_sel_is_5_o ;
  wire \picorv32_core/mux61_sel_is_5_o ;
  wire \picorv32_core/mux68_b0_sel_is_2_o ;
  wire \picorv32_core/mux69_b0_sel_is_1_o ;
  wire \picorv32_core/mux75_b0_sel_is_0_o ;
  wire \picorv32_core/mux76_b0_sel_is_2_o ;
  wire \picorv32_core/mux77_b0_sel_is_0_o ;
  wire \picorv32_core/mux77_b0_sel_is_0_o_neg ;
  wire \picorv32_core/mux77_b4_sel_is_2_o ;
  wire \picorv32_core/mux80_b0_sel_is_4_o ;
  wire \picorv32_core/mux80_b3_sel_is_4_o ;
  wire \picorv32_core/mux80_b4_sel_is_12_o ;
  wire \picorv32_core/mux81_sel_is_1_o ;
  wire \picorv32_core/mux84_sel_is_12_o ;
  wire \picorv32_core/mux88_b0_sel_is_2_o ;
  wire \picorv32_core/mux88_b0_sel_is_2_o_neg ;
  wire \picorv32_core/mux90_b1_sel_is_2_o ;
  wire \picorv32_core/mux90_b1_sel_is_2_o_neg ;
  wire \picorv32_core/mux91_b0_sel_is_0_o ;
  wire \picorv32_core/mux92_b1_sel_is_0_o ;
  wire \picorv32_core/mux93_b0_sel_is_2_o ;
  wire \picorv32_core/mux94_b0_sel_is_0_o ;
  wire \picorv32_core/n0 ;
  wire \picorv32_core/n1 ;
  wire \picorv32_core/n10 ;
  wire \picorv32_core/n100 ;
  wire \picorv32_core/n101 ;
  wire \picorv32_core/n104 ;
  wire \picorv32_core/n106 ;
  wire \picorv32_core/n11 ;
  wire \picorv32_core/n111 ;
  wire \picorv32_core/n111_neg ;
  wire \picorv32_core/n12 ;
  wire \picorv32_core/n120 ;
  wire \picorv32_core/n121 ;
  wire \picorv32_core/n125 ;
  wire \picorv32_core/n129 ;
  wire \picorv32_core/n13 ;
  wire \picorv32_core/n130 ;
  wire \picorv32_core/n131 ;
  wire \picorv32_core/n139 ;
  wire \picorv32_core/n14 ;
  wire \picorv32_core/n144 ;
  wire \picorv32_core/n148 ;
  wire \picorv32_core/n15 ;
  wire \picorv32_core/n16 ;
  wire \picorv32_core/n165 ;
  wire \picorv32_core/n166 ;
  wire \picorv32_core/n167 ;
  wire \picorv32_core/n168 ;
  wire \picorv32_core/n169 ;
  wire \picorv32_core/n170 ;
  wire \picorv32_core/n171 ;
  wire \picorv32_core/n172 ;
  wire \picorv32_core/n173 ;
  wire \picorv32_core/n174 ;
  wire \picorv32_core/n175 ;
  wire \picorv32_core/n176 ;
  wire \picorv32_core/n177 ;
  wire \picorv32_core/n178 ;
  wire \picorv32_core/n179 ;
  wire \picorv32_core/n18 ;
  wire \picorv32_core/n180 ;
  wire \picorv32_core/n181 ;
  wire \picorv32_core/n182 ;
  wire \picorv32_core/n183 ;
  wire \picorv32_core/n184 ;
  wire \picorv32_core/n185 ;
  wire \picorv32_core/n188 ;
  wire \picorv32_core/n19 ;
  wire \picorv32_core/n190 ;
  wire \picorv32_core/n191 ;
  wire \picorv32_core/n193 ;
  wire \picorv32_core/n193_neg ;
  wire \picorv32_core/n194 ;
  wire \picorv32_core/n197 ;
  wire \picorv32_core/n20 ;
  wire \picorv32_core/n201 ;
  wire \picorv32_core/n203 ;
  wire \picorv32_core/n203_neg ;
  wire \picorv32_core/n21 ;
  wire \picorv32_core/n211 ;
  wire \picorv32_core/n213 ;
  wire \picorv32_core/n22 ;
  wire \picorv32_core/n228 ;
  wire \picorv32_core/n233 ;
  wire \picorv32_core/n234 ;
  wire \picorv32_core/n238 ;
  wire \picorv32_core/n24 ;
  wire \picorv32_core/n240 ;
  wire \picorv32_core/n241 ;
  wire \picorv32_core/n249 ;
  wire \picorv32_core/n25 ;
  wire \picorv32_core/n250 ;
  wire \picorv32_core/n251 ;
  wire \picorv32_core/n252 ;
  wire \picorv32_core/n253 ;
  wire \picorv32_core/n254 ;
  wire \picorv32_core/n255 ;
  wire \picorv32_core/n256 ;
  wire \picorv32_core/n26 ;
  wire \picorv32_core/n273 ;
  wire \picorv32_core/n274 ;
  wire \picorv32_core/n274_neg ;
  wire \picorv32_core/n275 ;
  wire \picorv32_core/n276 ;
  wire \picorv32_core/n277 ;
  wire \picorv32_core/n278 ;
  wire \picorv32_core/n279 ;
  wire \picorv32_core/n28 ;
  wire \picorv32_core/n280 ;
  wire \picorv32_core/n281 ;
  wire \picorv32_core/n282 ;
  wire \picorv32_core/n283 ;
  wire \picorv32_core/n284 ;
  wire \picorv32_core/n285 ;
  wire \picorv32_core/n286 ;
  wire \picorv32_core/n287 ;
  wire \picorv32_core/n288 ;
  wire \picorv32_core/n289 ;
  wire \picorv32_core/n29 ;
  wire \picorv32_core/n290 ;
  wire \picorv32_core/n291 ;
  wire \picorv32_core/n292 ;
  wire \picorv32_core/n293 ;
  wire \picorv32_core/n294 ;
  wire \picorv32_core/n295 ;
  wire \picorv32_core/n296 ;
  wire \picorv32_core/n297 ;
  wire \picorv32_core/n298 ;
  wire \picorv32_core/n299 ;
  wire \picorv32_core/n300 ;
  wire \picorv32_core/n301 ;
  wire \picorv32_core/n302 ;
  wire \picorv32_core/n303 ;
  wire \picorv32_core/n304 ;
  wire \picorv32_core/n305 ;
  wire \picorv32_core/n306 ;
  wire \picorv32_core/n307 ;
  wire \picorv32_core/n308 ;
  wire \picorv32_core/n309 ;
  wire \picorv32_core/n310 ;
  wire \picorv32_core/n311 ;
  wire \picorv32_core/n312 ;
  wire \picorv32_core/n313 ;
  wire \picorv32_core/n314 ;
  wire \picorv32_core/n315 ;
  wire \picorv32_core/n316 ;
  wire \picorv32_core/n317 ;
  wire \picorv32_core/n318 ;
  wire \picorv32_core/n319 ;
  wire \picorv32_core/n320 ;
  wire \picorv32_core/n321 ;
  wire \picorv32_core/n322 ;
  wire \picorv32_core/n323 ;
  wire \picorv32_core/n324 ;
  wire \picorv32_core/n325 ;
  wire \picorv32_core/n326 ;
  wire \picorv32_core/n327 ;
  wire \picorv32_core/n328 ;
  wire \picorv32_core/n329 ;
  wire \picorv32_core/n330 ;
  wire \picorv32_core/n331 ;
  wire \picorv32_core/n332 ;
  wire \picorv32_core/n333 ;
  wire \picorv32_core/n334 ;
  wire \picorv32_core/n335 ;
  wire \picorv32_core/n336 ;
  wire \picorv32_core/n337 ;
  wire \picorv32_core/n338 ;
  wire \picorv32_core/n339 ;
  wire \picorv32_core/n340 ;
  wire \picorv32_core/n341 ;
  wire \picorv32_core/n342 ;
  wire \picorv32_core/n343 ;
  wire \picorv32_core/n344 ;
  wire \picorv32_core/n345 ;
  wire \picorv32_core/n346 ;
  wire \picorv32_core/n347 ;
  wire \picorv32_core/n348 ;
  wire \picorv32_core/n349 ;
  wire \picorv32_core/n350 ;
  wire \picorv32_core/n351 ;
  wire \picorv32_core/n353 ;
  wire \picorv32_core/n354 ;
  wire \picorv32_core/n356 ;
  wire \picorv32_core/n37 ;
  wire \picorv32_core/n4 ;
  wire \picorv32_core/n407 ;
  wire \picorv32_core/n43 ;
  wire \picorv32_core/n432 ;
  wire \picorv32_core/n436 ;
  wire \picorv32_core/n437 ;
  wire \picorv32_core/n438 ;
  wire \picorv32_core/n44 ;
  wire \picorv32_core/n440 ;
  wire \picorv32_core/n442 ;
  wire \picorv32_core/n444 ;
  wire \picorv32_core/n447 ;
  wire \picorv32_core/n448 ;
  wire \picorv32_core/n451 ;
  wire \picorv32_core/n452 ;
  wire \picorv32_core/n456 ;
  wire \picorv32_core/n457 ;
  wire \picorv32_core/n458 ;
  wire \picorv32_core/n46 ;
  wire \picorv32_core/n461 ;
  wire \picorv32_core/n462 ;
  wire \picorv32_core/n463 ;
  wire \picorv32_core/n464 ;
  wire \picorv32_core/n466 ;
  wire \picorv32_core/n467 ;
  wire \picorv32_core/n468 ;
  wire \picorv32_core/n469 ;
  wire \picorv32_core/n470 ;
  wire \picorv32_core/n471 ;
  wire \picorv32_core/n472 ;
  wire \picorv32_core/n473 ;
  wire \picorv32_core/n474 ;
  wire \picorv32_core/n475 ;
  wire \picorv32_core/n476 ;
  wire \picorv32_core/n477 ;
  wire \picorv32_core/n478 ;
  wire \picorv32_core/n479 ;
  wire \picorv32_core/n48 ;
  wire \picorv32_core/n480 ;
  wire \picorv32_core/n481 ;
  wire \picorv32_core/n482 ;
  wire \picorv32_core/n483 ;
  wire \picorv32_core/n484 ;
  wire \picorv32_core/n485 ;
  wire \picorv32_core/n486 ;
  wire \picorv32_core/n487 ;
  wire \picorv32_core/n488 ;
  wire \picorv32_core/n489 ;
  wire \picorv32_core/n490 ;
  wire \picorv32_core/n491 ;
  wire \picorv32_core/n492 ;
  wire \picorv32_core/n493 ;
  wire \picorv32_core/n494 ;
  wire \picorv32_core/n495 ;
  wire \picorv32_core/n497 ;
  wire \picorv32_core/n498 ;
  wire \picorv32_core/n499 ;
  wire \picorv32_core/n50 ;
  wire \picorv32_core/n505 ;
  wire \picorv32_core/n51 ;
  wire \picorv32_core/n513 ;
  wire \picorv32_core/n514 ;
  wire \picorv32_core/n519 ;
  wire \picorv32_core/n520 ;
  wire \picorv32_core/n522 ;
  wire \picorv32_core/n523 ;
  wire \picorv32_core/n526 ;
  wire \picorv32_core/n529 ;
  wire \picorv32_core/n530 ;
  wire \picorv32_core/n531 ;
  wire \picorv32_core/n533 ;
  wire \picorv32_core/n534 ;
  wire \picorv32_core/n535 ;
  wire \picorv32_core/n536 ;
  wire \picorv32_core/n537 ;
  wire \picorv32_core/n539 ;
  wire \picorv32_core/n54 ;
  wire \picorv32_core/n540 ;
  wire \picorv32_core/n541 ;
  wire \picorv32_core/n547 ;
  wire \picorv32_core/n548 ;
  wire \picorv32_core/n54_neg ;
  wire \picorv32_core/n550 ;
  wire \picorv32_core/n552 ;
  wire \picorv32_core/n553 ;
  wire \picorv32_core/n554 ;
  wire \picorv32_core/n555 ;
  wire \picorv32_core/n557 ;
  wire \picorv32_core/n56 ;
  wire \picorv32_core/n568 ;
  wire \picorv32_core/n56_neg ;
  wire \picorv32_core/n572 ;
  wire \picorv32_core/n573 ;
  wire \picorv32_core/n574 ;
  wire \picorv32_core/n58 ;
  wire \picorv32_core/n580 ;
  wire \picorv32_core/n588 ;
  wire \picorv32_core/n589 ;
  wire \picorv32_core/n58_neg ;
  wire \picorv32_core/n592 ;
  wire \picorv32_core/n593 ;
  wire \picorv32_core/n594 ;
  wire \picorv32_core/n595 ;
  wire \picorv32_core/n597 ;
  wire \picorv32_core/n598 ;
  wire \picorv32_core/n599 ;
  wire \picorv32_core/n600 ;
  wire \picorv32_core/n603 ;
  wire \picorv32_core/n605 ;
  wire \picorv32_core/n606 ;
  wire \picorv32_core/n607 ;
  wire \picorv32_core/n608 ;
  wire \picorv32_core/n609 ;
  wire \picorv32_core/n61 ;
  wire \picorv32_core/n610 ;
  wire \picorv32_core/n611 ;
  wire \picorv32_core/n612 ;
  wire \picorv32_core/n613 ;
  wire \picorv32_core/n614 ;
  wire \picorv32_core/n615 ;
  wire \picorv32_core/n616 ;
  wire \picorv32_core/n617 ;
  wire \picorv32_core/n618 ;
  wire \picorv32_core/n619 ;
  wire \picorv32_core/n61_neg ;
  wire \picorv32_core/n622 ;
  wire \picorv32_core/n623 ;
  wire \picorv32_core/n624 ;
  wire \picorv32_core/n625 ;
  wire \picorv32_core/n626 ;
  wire \picorv32_core/n627 ;
  wire \picorv32_core/n63 ;
  wire \picorv32_core/n632 ;
  wire \picorv32_core/n633 ;
  wire \picorv32_core/n639 ;
  wire \picorv32_core/n63_neg ;
  wire \picorv32_core/n640 ;
  wire \picorv32_core/n643 ;
  wire \picorv32_core/n644 ;
  wire \picorv32_core/n645 ;
  wire \picorv32_core/n646 ;
  wire \picorv32_core/n647 ;
  wire \picorv32_core/n648 ;
  wire \picorv32_core/n65 ;
  wire \picorv32_core/n650 ;
  wire \picorv32_core/n651 ;
  wire \picorv32_core/n653 ;
  wire \picorv32_core/n654 ;
  wire \picorv32_core/n655 ;
  wire \picorv32_core/n659 ;
  wire \picorv32_core/n65_neg ;
  wire \picorv32_core/n662 ;
  wire \picorv32_core/n663 ;
  wire \picorv32_core/n664 ;
  wire \picorv32_core/n665 ;
  wire \picorv32_core/n666 ;
  wire \picorv32_core/n667 ;
  wire \picorv32_core/n668 ;
  wire \picorv32_core/n669 ;
  wire \picorv32_core/n67 ;
  wire \picorv32_core/n670 ;
  wire \picorv32_core/n671 ;
  wire \picorv32_core/n675 ;
  wire \picorv32_core/n676 ;
  wire \picorv32_core/n677 ;
  wire \picorv32_core/n678 ;
  wire \picorv32_core/n679 ;
  wire \picorv32_core/n67_neg ;
  wire \picorv32_core/n680 ;
  wire \picorv32_core/n681 ;
  wire \picorv32_core/n682 ;
  wire \picorv32_core/n683 ;
  wire \picorv32_core/n684 ;
  wire \picorv32_core/n685 ;
  wire \picorv32_core/n686 ;
  wire \picorv32_core/n687 ;
  wire \picorv32_core/n697 ;
  wire \picorv32_core/n698 ;
  wire \picorv32_core/n7 ;
  wire \picorv32_core/n701 ;
  wire \picorv32_core/n701_neg ;
  wire \picorv32_core/n718 ;
  wire \picorv32_core/n72 ;
  wire \picorv32_core/n727 ;
  wire \picorv32_core/n728 ;
  wire \picorv32_core/n729 ;
  wire \picorv32_core/n73 ;
  wire \picorv32_core/n731 ;
  wire \picorv32_core/n732 ;
  wire \picorv32_core/n733 ;
  wire \picorv32_core/n734 ;
  wire \picorv32_core/n735 ;
  wire \picorv32_core/n736 ;
  wire \picorv32_core/n736_neg ;
  wire \picorv32_core/n738 ;
  wire \picorv32_core/n739 ;
  wire \picorv32_core/n74 ;
  wire \picorv32_core/n740 ;
  wire \picorv32_core/n740_neg ;
  wire \picorv32_core/n743 ;
  wire \picorv32_core/n744 ;
  wire \picorv32_core/n744_neg ;
  wire \picorv32_core/n746 ;
  wire \picorv32_core/n747 ;
  wire \picorv32_core/n749 ;
  wire \picorv32_core/n74_neg ;
  wire \picorv32_core/n79 ;
  wire \picorv32_core/n8 ;
  wire \picorv32_core/n80 ;
  wire \picorv32_core/n80_neg ;
  wire \picorv32_core/n84 ;
  wire \picorv32_core/n85 ;
  wire \picorv32_core/n86 ;
  wire \picorv32_core/n87 ;
  wire \picorv32_core/n87_neg ;
  wire \picorv32_core/n9 ;
  wire \picorv32_core/n92 ;
  wire \picorv32_core/n92_neg ;
  wire \picorv32_core/n96 ;
  wire \picorv32_core/n97 ;
  wire \picorv32_core/n98 ;
  wire \picorv32_core/n99 ;
  wire \picorv32_core/pcpi_rs1$0$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$1$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$10$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$11$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$12$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$13$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$14$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$15$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$16$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$17$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$18$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$19$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$2$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$20$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$21$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$22$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$23$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$24$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$25$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$26$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$27$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$28$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$29$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$3$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$30$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$31$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$4$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$5$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$6$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$7$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$8$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs1$9$ ;  // ../src/picorv32.v(96)
  wire \picorv32_core/pcpi_rs2$10$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$11$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$12$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$13$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$14$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$15$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$16$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$17$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$18$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$19$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$20$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$21$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$22$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$23$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$24$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$25$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$26$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$27$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$28$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$29$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$30$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$31$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$8$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/pcpi_rs2$9$ ;  // ../src/picorv32.v(97)
  wire \picorv32_core/prefetched_high_word ;  // ../src/picorv32.v(329)
  wire \picorv32_core/sel11_b1/or_B1_B2_o ;
  wire \picorv32_core/sel11_b1/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b10/or_B1_B2_o ;
  wire \picorv32_core/sel11_b10/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b11/or_B1_B2_o ;
  wire \picorv32_core/sel11_b11/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b12/or_B1_B2_o ;
  wire \picorv32_core/sel11_b12/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b12/or_B4_B5_o ;
  wire \picorv32_core/sel11_b13/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b13/or_B4_B5_o ;
  wire \picorv32_core/sel11_b14/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b14/or_B4_B5_o ;
  wire \picorv32_core/sel11_b15/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b15/or_B4_B5_o ;
  wire \picorv32_core/sel11_b16/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b16/or_B4_B5_o ;
  wire \picorv32_core/sel11_b17/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b17/or_B4_B5_o ;
  wire \picorv32_core/sel11_b18/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b18/or_B4_B5_o ;
  wire \picorv32_core/sel11_b19/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b19/or_B4_B5_o ;
  wire \picorv32_core/sel11_b2/or_B1_B2_o ;
  wire \picorv32_core/sel11_b2/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b20/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b20/or_B4_B5_o ;
  wire \picorv32_core/sel11_b21/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b21/or_B4_B5_o ;
  wire \picorv32_core/sel11_b22/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b22/or_B4_B5_o ;
  wire \picorv32_core/sel11_b23/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b23/or_B4_B5_o ;
  wire \picorv32_core/sel11_b24/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b24/or_B4_B5_o ;
  wire \picorv32_core/sel11_b25/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b25/or_B4_B5_o ;
  wire \picorv32_core/sel11_b26/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b26/or_B4_B5_o ;
  wire \picorv32_core/sel11_b27/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b27/or_B4_B5_o ;
  wire \picorv32_core/sel11_b28/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b28/or_B4_B5_o ;
  wire \picorv32_core/sel11_b29/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b29/or_B4_B5_o ;
  wire \picorv32_core/sel11_b3/or_B1_B2_o ;
  wire \picorv32_core/sel11_b3/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b30/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b30/or_B4_B5_o ;
  wire \picorv32_core/sel11_b31/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b31/or_B4_B5_o ;
  wire \picorv32_core/sel11_b4/or_B1_B2_o ;
  wire \picorv32_core/sel11_b4/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b5/or_B1_B2_o ;
  wire \picorv32_core/sel11_b5/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b6/or_B1_B2_o ;
  wire \picorv32_core/sel11_b6/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b7/or_B1_B2_o ;
  wire \picorv32_core/sel11_b7/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b8/or_B1_B2_o ;
  wire \picorv32_core/sel11_b8/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel11_b9/or_B1_B2_o ;
  wire \picorv32_core/sel11_b9/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel12/or_B0_or_B1_B2_o_o ;
  wire \picorv32_core/sel12/or_B1_B2_o ;
  wire \picorv32_core/sel12/or_B3_or_B4_B5_o_o ;
  wire \picorv32_core/sel12/or_B4_B5_o ;
  wire \picorv32_core/sel13_b0/or_B0_B1_o ;
  wire \picorv32_core/sel13_b0/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b0/or_B3_B4_o ;
  wire \picorv32_core/sel13_b1/or_B0_B1_o ;
  wire \picorv32_core/sel13_b1/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b10/or_B0_B1_o ;
  wire \picorv32_core/sel13_b10/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b11/or_B0_B1_o ;
  wire \picorv32_core/sel13_b11/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b12/or_B0_B1_o ;
  wire \picorv32_core/sel13_b12/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b13/or_B0_B1_o ;
  wire \picorv32_core/sel13_b13/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b14/or_B0_B1_o ;
  wire \picorv32_core/sel13_b14/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b15/or_B0_B1_o ;
  wire \picorv32_core/sel13_b15/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b16/or_B0_B1_o ;
  wire \picorv32_core/sel13_b16/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b17/or_B0_B1_o ;
  wire \picorv32_core/sel13_b17/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b18/or_B0_B1_o ;
  wire \picorv32_core/sel13_b18/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b19/or_B0_B1_o ;
  wire \picorv32_core/sel13_b19/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b2/or_B0_B1_o ;
  wire \picorv32_core/sel13_b2/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b20/or_B0_B1_o ;
  wire \picorv32_core/sel13_b20/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b21/or_B0_B1_o ;
  wire \picorv32_core/sel13_b21/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b22/or_B0_B1_o ;
  wire \picorv32_core/sel13_b22/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b23/or_B0_B1_o ;
  wire \picorv32_core/sel13_b23/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b24/or_B0_B1_o ;
  wire \picorv32_core/sel13_b24/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b25/or_B0_B1_o ;
  wire \picorv32_core/sel13_b25/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b26/or_B0_B1_o ;
  wire \picorv32_core/sel13_b26/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b27/or_B0_B1_o ;
  wire \picorv32_core/sel13_b27/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b28/or_B0_B1_o ;
  wire \picorv32_core/sel13_b28/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b29/or_B0_B1_o ;
  wire \picorv32_core/sel13_b29/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b3/or_B0_B1_o ;
  wire \picorv32_core/sel13_b3/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b30/or_B0_B1_o ;
  wire \picorv32_core/sel13_b30/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b31/or_B0_B1_o ;
  wire \picorv32_core/sel13_b31/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b4/or_B0_B1_o ;
  wire \picorv32_core/sel13_b4/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b5/or_B0_B1_o ;
  wire \picorv32_core/sel13_b5/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b6/or_B0_B1_o ;
  wire \picorv32_core/sel13_b6/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b7/or_B0_B1_o ;
  wire \picorv32_core/sel13_b7/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b8/or_B0_B1_o ;
  wire \picorv32_core/sel13_b8/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel13_b9/or_B0_B1_o ;
  wire \picorv32_core/sel13_b9/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel15_b0_sel_is_3_o ;
  wire \picorv32_core/sel16_b0/or_B0_B1_o ;
  wire \picorv32_core/sel16_b0/or_B2_B3_o ;
  wire \picorv32_core/sel16_b1/or_B0_B1_o ;
  wire \picorv32_core/sel16_b1/or_B2_B3_o ;
  wire \picorv32_core/sel16_b10/or_B0_B1_o ;
  wire \picorv32_core/sel16_b10/or_B2_B3_o ;
  wire \picorv32_core/sel16_b11/or_B0_B1_o ;
  wire \picorv32_core/sel16_b11/or_B2_B3_o ;
  wire \picorv32_core/sel16_b12/or_B0_B1_o ;
  wire \picorv32_core/sel16_b12/or_B2_B3_o ;
  wire \picorv32_core/sel16_b13/or_B0_B1_o ;
  wire \picorv32_core/sel16_b13/or_B2_B3_o ;
  wire \picorv32_core/sel16_b14/or_B0_B1_o ;
  wire \picorv32_core/sel16_b14/or_B2_B3_o ;
  wire \picorv32_core/sel16_b15/or_B0_B1_o ;
  wire \picorv32_core/sel16_b15/or_B2_B3_o ;
  wire \picorv32_core/sel16_b16/or_B0_B1_o ;
  wire \picorv32_core/sel16_b16/or_B2_B3_o ;
  wire \picorv32_core/sel16_b17/or_B0_B1_o ;
  wire \picorv32_core/sel16_b17/or_B2_B3_o ;
  wire \picorv32_core/sel16_b18/or_B0_B1_o ;
  wire \picorv32_core/sel16_b18/or_B2_B3_o ;
  wire \picorv32_core/sel16_b19/or_B0_B1_o ;
  wire \picorv32_core/sel16_b19/or_B2_B3_o ;
  wire \picorv32_core/sel16_b2/or_B0_B1_o ;
  wire \picorv32_core/sel16_b2/or_B2_B3_o ;
  wire \picorv32_core/sel16_b20/or_B0_B1_o ;
  wire \picorv32_core/sel16_b20/or_B2_B3_o ;
  wire \picorv32_core/sel16_b21/or_B0_B1_o ;
  wire \picorv32_core/sel16_b21/or_B2_B3_o ;
  wire \picorv32_core/sel16_b22/or_B0_B1_o ;
  wire \picorv32_core/sel16_b22/or_B2_B3_o ;
  wire \picorv32_core/sel16_b23/or_B0_B1_o ;
  wire \picorv32_core/sel16_b23/or_B2_B3_o ;
  wire \picorv32_core/sel16_b24/or_B0_B1_o ;
  wire \picorv32_core/sel16_b24/or_B2_B3_o ;
  wire \picorv32_core/sel16_b25/or_B0_B1_o ;
  wire \picorv32_core/sel16_b25/or_B2_B3_o ;
  wire \picorv32_core/sel16_b26/or_B0_B1_o ;
  wire \picorv32_core/sel16_b26/or_B2_B3_o ;
  wire \picorv32_core/sel16_b27/or_B0_B1_o ;
  wire \picorv32_core/sel16_b27/or_B2_B3_o ;
  wire \picorv32_core/sel16_b28/or_B0_B1_o ;
  wire \picorv32_core/sel16_b28/or_B2_B3_o ;
  wire \picorv32_core/sel16_b29/or_B0_B1_o ;
  wire \picorv32_core/sel16_b29/or_B2_B3_o ;
  wire \picorv32_core/sel16_b3/or_B0_B1_o ;
  wire \picorv32_core/sel16_b3/or_B2_B3_o ;
  wire \picorv32_core/sel16_b30/or_B0_B1_o ;
  wire \picorv32_core/sel16_b30/or_B2_B3_o ;
  wire \picorv32_core/sel16_b31/or_B0_B1_o ;
  wire \picorv32_core/sel16_b31/or_B2_B3_o ;
  wire \picorv32_core/sel16_b4/or_B0_B1_o ;
  wire \picorv32_core/sel16_b4/or_B2_B3_o ;
  wire \picorv32_core/sel16_b5/or_B0_B1_o ;
  wire \picorv32_core/sel16_b5/or_B2_B3_o ;
  wire \picorv32_core/sel16_b6/or_B0_B1_o ;
  wire \picorv32_core/sel16_b6/or_B2_B3_o ;
  wire \picorv32_core/sel16_b7/or_B0_B1_o ;
  wire \picorv32_core/sel16_b7/or_B2_B3_o ;
  wire \picorv32_core/sel16_b8/or_B0_B1_o ;
  wire \picorv32_core/sel16_b8/or_B2_B3_o ;
  wire \picorv32_core/sel16_b9/or_B0_B1_o ;
  wire \picorv32_core/sel16_b9/or_B2_B3_o ;
  wire \picorv32_core/sel18/or_B1_B2_o ;
  wire \picorv32_core/sel19_b2/or_B0_or_B1_B2_o_o ;
  wire \picorv32_core/sel19_b3/or_B0_or_B1_B2_o_o ;
  wire \picorv32_core/sel2/or_B1_B2_o ;
  wire \picorv32_core/sel23/or_B0_B1_o ;
  wire \picorv32_core/sel23/or_B2_B3_o ;
  wire \picorv32_core/sel27_b16/or_B1_B2_o ;
  wire \picorv32_core/sel27_b17/or_B1_B2_o ;
  wire \picorv32_core/sel27_b18/or_B1_B2_o ;
  wire \picorv32_core/sel27_b19/or_B1_B2_o ;
  wire \picorv32_core/sel27_b20/or_B1_B2_o ;
  wire \picorv32_core/sel27_b21/or_B1_B2_o ;
  wire \picorv32_core/sel27_b22/or_B1_B2_o ;
  wire \picorv32_core/sel27_b23/or_B1_B2_o ;
  wire \picorv32_core/sel27_b24/or_B1_B2_o ;
  wire \picorv32_core/sel27_b25/or_B1_B2_o ;
  wire \picorv32_core/sel27_b26/or_B1_B2_o ;
  wire \picorv32_core/sel27_b27/or_B1_B2_o ;
  wire \picorv32_core/sel27_b28/or_B1_B2_o ;
  wire \picorv32_core/sel27_b29/or_B1_B2_o ;
  wire \picorv32_core/sel27_b30/or_B1_B2_o ;
  wire \picorv32_core/sel27_b31/or_B1_B2_o ;
  wire \picorv32_core/sel28/or_B0_B1_o ;
  wire \picorv32_core/sel28/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel28/or_B3_B4_o ;
  wire \picorv32_core/sel29_b0/or_B0_B1_o ;
  wire \picorv32_core/sel29_b0/or_B2_B3_o ;
  wire \picorv32_core/sel29_b0/or_B4_B5_o ;
  wire \picorv32_core/sel29_b0/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel29_b0/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel29_b1/or_B0_B1_o ;
  wire \picorv32_core/sel29_b1/or_B2_B3_o ;
  wire \picorv32_core/sel29_b1/or_B4_B5_o ;
  wire \picorv32_core/sel29_b1/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel29_b1/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel32/or_B0_B1_o ;
  wire \picorv32_core/sel32/or_B2_or_B3_B4_o_o ;
  wire \picorv32_core/sel34/or_B1_B2_o ;
  wire \picorv32_core/sel38_b0/or_B0_B1_o ;
  wire \picorv32_core/sel38_b0/or_B2_B3_o ;
  wire \picorv32_core/sel38_b0/or_B4_B5_o ;
  wire \picorv32_core/sel38_b0/or_B6_B7_o ;
  wire \picorv32_core/sel38_b0/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel38_b0/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel38_b1/or_B0_B1_o ;
  wire \picorv32_core/sel38_b1/or_B2_B3_o ;
  wire \picorv32_core/sel38_b1/or_B4_B5_o ;
  wire \picorv32_core/sel38_b1/or_B6_B7_o ;
  wire \picorv32_core/sel38_b1/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel38_b1/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel38_b2/or_B0_B1_o ;
  wire \picorv32_core/sel38_b2/or_B2_B3_o ;
  wire \picorv32_core/sel38_b2/or_B4_B5_o ;
  wire \picorv32_core/sel38_b2/or_B6_B7_o ;
  wire \picorv32_core/sel38_b2/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel38_b2/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel38_b3/or_B0_B1_o ;
  wire \picorv32_core/sel38_b3/or_B2_B3_o ;
  wire \picorv32_core/sel38_b3/or_B4_B5_o ;
  wire \picorv32_core/sel38_b3/or_B6_B7_o ;
  wire \picorv32_core/sel38_b3/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel38_b3/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel38_b4/or_B0_B1_o ;
  wire \picorv32_core/sel38_b4/or_B2_B3_o ;
  wire \picorv32_core/sel38_b4/or_B4_B5_o ;
  wire \picorv32_core/sel38_b4/or_B6_B7_o ;
  wire \picorv32_core/sel38_b4/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel38_b4/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel39_b0_sel_is_3_o ;
  wire \picorv32_core/sel40_b0/or_B0_B1_o ;
  wire \picorv32_core/sel40_b0/or_B2_B3_o ;
  wire \picorv32_core/sel40_b0/or_B6_B7_o ;
  wire \picorv32_core/sel40_b0/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel40_b0/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel40_b1/or_B0_B1_o ;
  wire \picorv32_core/sel40_b1/or_B2_B3_o ;
  wire \picorv32_core/sel40_b1/or_B4_B5_o ;
  wire \picorv32_core/sel40_b1/or_B6_B7_o ;
  wire \picorv32_core/sel40_b1/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel40_b1/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel40_b2/or_B0_B1_o ;
  wire \picorv32_core/sel40_b2/or_B2_B3_o ;
  wire \picorv32_core/sel40_b2/or_B4_B5_o ;
  wire \picorv32_core/sel40_b2/or_B6_B7_o ;
  wire \picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel40_b2/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel40_b3/or_B0_B1_o ;
  wire \picorv32_core/sel40_b3/or_B2_B3_o ;
  wire \picorv32_core/sel40_b3/or_B4_B5_o ;
  wire \picorv32_core/sel40_b3/or_B6_B7_o ;
  wire \picorv32_core/sel40_b3/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel40_b3/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel40_b4/or_B0_B1_o ;
  wire \picorv32_core/sel40_b4/or_B2_B3_o ;
  wire \picorv32_core/sel40_b4/or_B6_B7_o ;
  wire \picorv32_core/sel40_b4/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel40_b5/or_B0_B1_o ;
  wire \picorv32_core/sel40_b5/or_B2_B3_o ;
  wire \picorv32_core/sel40_b5/or_B6_B7_o ;
  wire \picorv32_core/sel40_b5/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel40_b6/or_B0_B1_o ;
  wire \picorv32_core/sel40_b6/or_B2_B3_o ;
  wire \picorv32_core/sel40_b6/or_B6_B7_o ;
  wire \picorv32_core/sel40_b6/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel40_b6/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel40_b7/or_B0_B1_o ;
  wire \picorv32_core/sel40_b7/or_B2_B3_o ;
  wire \picorv32_core/sel40_b7/or_B6_B7_o ;
  wire \picorv32_core/sel40_b7/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel40_b7/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b0/or_B0_B1_o ;
  wire \picorv32_core/sel41_b0/or_B2_B3_o ;
  wire \picorv32_core/sel41_b0/or_B4_B5_o ;
  wire \picorv32_core/sel41_b0/or_B6_B7_o ;
  wire \picorv32_core/sel41_b0/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b0/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b1/or_B0_B1_o ;
  wire \picorv32_core/sel41_b1/or_B2_B3_o ;
  wire \picorv32_core/sel41_b1/or_B4_B5_o ;
  wire \picorv32_core/sel41_b1/or_B6_B7_o ;
  wire \picorv32_core/sel41_b1/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b1/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b10/or_B0_B1_o ;
  wire \picorv32_core/sel41_b10/or_B2_B3_o ;
  wire \picorv32_core/sel41_b10/or_B4_B5_o ;
  wire \picorv32_core/sel41_b10/or_B6_B7_o ;
  wire \picorv32_core/sel41_b10/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b10/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b11/or_B0_B1_o ;
  wire \picorv32_core/sel41_b11/or_B2_B3_o ;
  wire \picorv32_core/sel41_b11/or_B4_B5_o ;
  wire \picorv32_core/sel41_b11/or_B6_B7_o ;
  wire \picorv32_core/sel41_b11/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b11/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b12/or_B0_B1_o ;
  wire \picorv32_core/sel41_b12/or_B2_B3_o ;
  wire \picorv32_core/sel41_b12/or_B4_B5_o ;
  wire \picorv32_core/sel41_b12/or_B6_B7_o ;
  wire \picorv32_core/sel41_b12/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b12/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b13/or_B0_B1_o ;
  wire \picorv32_core/sel41_b13/or_B2_B3_o ;
  wire \picorv32_core/sel41_b13/or_B4_B5_o ;
  wire \picorv32_core/sel41_b13/or_B6_B7_o ;
  wire \picorv32_core/sel41_b13/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b13/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b14/or_B0_B1_o ;
  wire \picorv32_core/sel41_b14/or_B2_B3_o ;
  wire \picorv32_core/sel41_b14/or_B4_B5_o ;
  wire \picorv32_core/sel41_b14/or_B6_B7_o ;
  wire \picorv32_core/sel41_b14/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b14/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b15/or_B0_B1_o ;
  wire \picorv32_core/sel41_b15/or_B2_B3_o ;
  wire \picorv32_core/sel41_b15/or_B4_B5_o ;
  wire \picorv32_core/sel41_b15/or_B6_B7_o ;
  wire \picorv32_core/sel41_b15/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b15/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b16/or_B0_B1_o ;
  wire \picorv32_core/sel41_b16/or_B2_B3_o ;
  wire \picorv32_core/sel41_b16/or_B4_B5_o ;
  wire \picorv32_core/sel41_b16/or_B6_B7_o ;
  wire \picorv32_core/sel41_b16/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b16/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b17/or_B0_B1_o ;
  wire \picorv32_core/sel41_b17/or_B2_B3_o ;
  wire \picorv32_core/sel41_b17/or_B4_B5_o ;
  wire \picorv32_core/sel41_b17/or_B6_B7_o ;
  wire \picorv32_core/sel41_b17/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b17/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b18/or_B0_B1_o ;
  wire \picorv32_core/sel41_b18/or_B2_B3_o ;
  wire \picorv32_core/sel41_b18/or_B4_B5_o ;
  wire \picorv32_core/sel41_b18/or_B6_B7_o ;
  wire \picorv32_core/sel41_b18/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b18/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b19/or_B0_B1_o ;
  wire \picorv32_core/sel41_b19/or_B2_B3_o ;
  wire \picorv32_core/sel41_b19/or_B4_B5_o ;
  wire \picorv32_core/sel41_b19/or_B6_B7_o ;
  wire \picorv32_core/sel41_b19/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b19/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b2/or_B0_B1_o ;
  wire \picorv32_core/sel41_b2/or_B2_B3_o ;
  wire \picorv32_core/sel41_b2/or_B4_B5_o ;
  wire \picorv32_core/sel41_b2/or_B6_B7_o ;
  wire \picorv32_core/sel41_b2/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b2/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b20/or_B0_B1_o ;
  wire \picorv32_core/sel41_b20/or_B2_B3_o ;
  wire \picorv32_core/sel41_b20/or_B4_B5_o ;
  wire \picorv32_core/sel41_b20/or_B6_B7_o ;
  wire \picorv32_core/sel41_b20/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b20/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b21/or_B0_B1_o ;
  wire \picorv32_core/sel41_b21/or_B2_B3_o ;
  wire \picorv32_core/sel41_b21/or_B4_B5_o ;
  wire \picorv32_core/sel41_b21/or_B6_B7_o ;
  wire \picorv32_core/sel41_b21/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b21/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b22/or_B0_B1_o ;
  wire \picorv32_core/sel41_b22/or_B2_B3_o ;
  wire \picorv32_core/sel41_b22/or_B4_B5_o ;
  wire \picorv32_core/sel41_b22/or_B6_B7_o ;
  wire \picorv32_core/sel41_b22/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b22/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b23/or_B0_B1_o ;
  wire \picorv32_core/sel41_b23/or_B2_B3_o ;
  wire \picorv32_core/sel41_b23/or_B4_B5_o ;
  wire \picorv32_core/sel41_b23/or_B6_B7_o ;
  wire \picorv32_core/sel41_b23/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b23/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b24/or_B0_B1_o ;
  wire \picorv32_core/sel41_b24/or_B2_B3_o ;
  wire \picorv32_core/sel41_b24/or_B4_B5_o ;
  wire \picorv32_core/sel41_b24/or_B6_B7_o ;
  wire \picorv32_core/sel41_b24/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b24/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b25/or_B0_B1_o ;
  wire \picorv32_core/sel41_b25/or_B2_B3_o ;
  wire \picorv32_core/sel41_b25/or_B4_B5_o ;
  wire \picorv32_core/sel41_b25/or_B6_B7_o ;
  wire \picorv32_core/sel41_b25/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b25/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b26/or_B0_B1_o ;
  wire \picorv32_core/sel41_b26/or_B2_B3_o ;
  wire \picorv32_core/sel41_b26/or_B4_B5_o ;
  wire \picorv32_core/sel41_b26/or_B6_B7_o ;
  wire \picorv32_core/sel41_b26/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b26/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b27/or_B0_B1_o ;
  wire \picorv32_core/sel41_b27/or_B2_B3_o ;
  wire \picorv32_core/sel41_b27/or_B4_B5_o ;
  wire \picorv32_core/sel41_b27/or_B6_B7_o ;
  wire \picorv32_core/sel41_b27/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b27/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b28/or_B0_B1_o ;
  wire \picorv32_core/sel41_b28/or_B2_B3_o ;
  wire \picorv32_core/sel41_b28/or_B4_B5_o ;
  wire \picorv32_core/sel41_b28/or_B6_B7_o ;
  wire \picorv32_core/sel41_b28/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b28/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b29/or_B0_B1_o ;
  wire \picorv32_core/sel41_b29/or_B2_B3_o ;
  wire \picorv32_core/sel41_b29/or_B4_B5_o ;
  wire \picorv32_core/sel41_b29/or_B6_B7_o ;
  wire \picorv32_core/sel41_b29/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b29/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b3/or_B0_B1_o ;
  wire \picorv32_core/sel41_b3/or_B2_B3_o ;
  wire \picorv32_core/sel41_b3/or_B4_B5_o ;
  wire \picorv32_core/sel41_b3/or_B6_B7_o ;
  wire \picorv32_core/sel41_b3/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b3/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b30/or_B0_B1_o ;
  wire \picorv32_core/sel41_b30/or_B2_B3_o ;
  wire \picorv32_core/sel41_b30/or_B4_B5_o ;
  wire \picorv32_core/sel41_b30/or_B6_B7_o ;
  wire \picorv32_core/sel41_b30/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b30/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b31/or_B0_B1_o ;
  wire \picorv32_core/sel41_b31/or_B2_B3_o ;
  wire \picorv32_core/sel41_b31/or_B4_B5_o ;
  wire \picorv32_core/sel41_b31/or_B6_B7_o ;
  wire \picorv32_core/sel41_b31/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b31/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b4/or_B0_B1_o ;
  wire \picorv32_core/sel41_b4/or_B2_B3_o ;
  wire \picorv32_core/sel41_b4/or_B4_B5_o ;
  wire \picorv32_core/sel41_b4/or_B6_B7_o ;
  wire \picorv32_core/sel41_b4/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b4/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b5/or_B0_B1_o ;
  wire \picorv32_core/sel41_b5/or_B2_B3_o ;
  wire \picorv32_core/sel41_b5/or_B4_B5_o ;
  wire \picorv32_core/sel41_b5/or_B6_B7_o ;
  wire \picorv32_core/sel41_b5/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b5/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b6/or_B0_B1_o ;
  wire \picorv32_core/sel41_b6/or_B2_B3_o ;
  wire \picorv32_core/sel41_b6/or_B4_B5_o ;
  wire \picorv32_core/sel41_b6/or_B6_B7_o ;
  wire \picorv32_core/sel41_b6/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b6/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b7/or_B0_B1_o ;
  wire \picorv32_core/sel41_b7/or_B2_B3_o ;
  wire \picorv32_core/sel41_b7/or_B4_B5_o ;
  wire \picorv32_core/sel41_b7/or_B6_B7_o ;
  wire \picorv32_core/sel41_b7/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b7/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b8/or_B0_B1_o ;
  wire \picorv32_core/sel41_b8/or_B2_B3_o ;
  wire \picorv32_core/sel41_b8/or_B4_B5_o ;
  wire \picorv32_core/sel41_b8/or_B6_B7_o ;
  wire \picorv32_core/sel41_b8/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b8/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel41_b9/or_B0_B1_o ;
  wire \picorv32_core/sel41_b9/or_B2_B3_o ;
  wire \picorv32_core/sel41_b9/or_B4_B5_o ;
  wire \picorv32_core/sel41_b9/or_B6_B7_o ;
  wire \picorv32_core/sel41_b9/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel41_b9/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b0/or_B0_B1_o ;
  wire \picorv32_core/sel42_b0/or_B2_B3_o ;
  wire \picorv32_core/sel42_b0/or_B4_B5_o ;
  wire \picorv32_core/sel42_b0/or_B6_B7_o ;
  wire \picorv32_core/sel42_b0/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b0/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b1/or_B0_B1_o ;
  wire \picorv32_core/sel42_b1/or_B2_B3_o ;
  wire \picorv32_core/sel42_b1/or_B4_B5_o ;
  wire \picorv32_core/sel42_b1/or_B6_B7_o ;
  wire \picorv32_core/sel42_b1/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b1/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b10/or_B0_B1_o ;
  wire \picorv32_core/sel42_b10/or_B2_B3_o ;
  wire \picorv32_core/sel42_b10/or_B4_B5_o ;
  wire \picorv32_core/sel42_b10/or_B6_B7_o ;
  wire \picorv32_core/sel42_b10/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b10/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b11/or_B0_B1_o ;
  wire \picorv32_core/sel42_b11/or_B2_B3_o ;
  wire \picorv32_core/sel42_b11/or_B4_B5_o ;
  wire \picorv32_core/sel42_b11/or_B6_B7_o ;
  wire \picorv32_core/sel42_b11/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b11/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b12/or_B0_B1_o ;
  wire \picorv32_core/sel42_b12/or_B2_B3_o ;
  wire \picorv32_core/sel42_b12/or_B4_B5_o ;
  wire \picorv32_core/sel42_b12/or_B6_B7_o ;
  wire \picorv32_core/sel42_b12/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b12/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b13/or_B0_B1_o ;
  wire \picorv32_core/sel42_b13/or_B2_B3_o ;
  wire \picorv32_core/sel42_b13/or_B4_B5_o ;
  wire \picorv32_core/sel42_b13/or_B6_B7_o ;
  wire \picorv32_core/sel42_b13/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b13/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b14/or_B0_B1_o ;
  wire \picorv32_core/sel42_b14/or_B2_B3_o ;
  wire \picorv32_core/sel42_b14/or_B4_B5_o ;
  wire \picorv32_core/sel42_b14/or_B6_B7_o ;
  wire \picorv32_core/sel42_b14/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b14/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b15/or_B0_B1_o ;
  wire \picorv32_core/sel42_b15/or_B2_B3_o ;
  wire \picorv32_core/sel42_b15/or_B4_B5_o ;
  wire \picorv32_core/sel42_b15/or_B6_B7_o ;
  wire \picorv32_core/sel42_b15/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b15/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b16/or_B0_B1_o ;
  wire \picorv32_core/sel42_b16/or_B2_B3_o ;
  wire \picorv32_core/sel42_b16/or_B4_B5_o ;
  wire \picorv32_core/sel42_b16/or_B6_B7_o ;
  wire \picorv32_core/sel42_b16/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b16/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b17/or_B0_B1_o ;
  wire \picorv32_core/sel42_b17/or_B2_B3_o ;
  wire \picorv32_core/sel42_b17/or_B4_B5_o ;
  wire \picorv32_core/sel42_b17/or_B6_B7_o ;
  wire \picorv32_core/sel42_b17/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b17/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b18/or_B0_B1_o ;
  wire \picorv32_core/sel42_b18/or_B2_B3_o ;
  wire \picorv32_core/sel42_b18/or_B4_B5_o ;
  wire \picorv32_core/sel42_b18/or_B6_B7_o ;
  wire \picorv32_core/sel42_b18/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b18/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b19/or_B0_B1_o ;
  wire \picorv32_core/sel42_b19/or_B2_B3_o ;
  wire \picorv32_core/sel42_b19/or_B4_B5_o ;
  wire \picorv32_core/sel42_b19/or_B6_B7_o ;
  wire \picorv32_core/sel42_b19/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b19/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b2/or_B0_B1_o ;
  wire \picorv32_core/sel42_b2/or_B2_B3_o ;
  wire \picorv32_core/sel42_b2/or_B4_B5_o ;
  wire \picorv32_core/sel42_b2/or_B6_B7_o ;
  wire \picorv32_core/sel42_b2/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b2/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b20/or_B0_B1_o ;
  wire \picorv32_core/sel42_b20/or_B2_B3_o ;
  wire \picorv32_core/sel42_b20/or_B4_B5_o ;
  wire \picorv32_core/sel42_b20/or_B6_B7_o ;
  wire \picorv32_core/sel42_b20/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b20/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b21/or_B0_B1_o ;
  wire \picorv32_core/sel42_b21/or_B2_B3_o ;
  wire \picorv32_core/sel42_b21/or_B4_B5_o ;
  wire \picorv32_core/sel42_b21/or_B6_B7_o ;
  wire \picorv32_core/sel42_b21/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b21/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b22/or_B0_B1_o ;
  wire \picorv32_core/sel42_b22/or_B2_B3_o ;
  wire \picorv32_core/sel42_b22/or_B4_B5_o ;
  wire \picorv32_core/sel42_b22/or_B6_B7_o ;
  wire \picorv32_core/sel42_b22/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b22/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b23/or_B0_B1_o ;
  wire \picorv32_core/sel42_b23/or_B2_B3_o ;
  wire \picorv32_core/sel42_b23/or_B4_B5_o ;
  wire \picorv32_core/sel42_b23/or_B6_B7_o ;
  wire \picorv32_core/sel42_b23/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b23/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b24/or_B0_B1_o ;
  wire \picorv32_core/sel42_b24/or_B2_B3_o ;
  wire \picorv32_core/sel42_b24/or_B4_B5_o ;
  wire \picorv32_core/sel42_b24/or_B6_B7_o ;
  wire \picorv32_core/sel42_b24/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b24/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b25/or_B0_B1_o ;
  wire \picorv32_core/sel42_b25/or_B2_B3_o ;
  wire \picorv32_core/sel42_b25/or_B4_B5_o ;
  wire \picorv32_core/sel42_b25/or_B6_B7_o ;
  wire \picorv32_core/sel42_b25/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b25/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b26/or_B0_B1_o ;
  wire \picorv32_core/sel42_b26/or_B2_B3_o ;
  wire \picorv32_core/sel42_b26/or_B4_B5_o ;
  wire \picorv32_core/sel42_b26/or_B6_B7_o ;
  wire \picorv32_core/sel42_b26/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b26/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b27/or_B0_B1_o ;
  wire \picorv32_core/sel42_b27/or_B2_B3_o ;
  wire \picorv32_core/sel42_b27/or_B4_B5_o ;
  wire \picorv32_core/sel42_b27/or_B6_B7_o ;
  wire \picorv32_core/sel42_b27/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b27/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b28/or_B0_B1_o ;
  wire \picorv32_core/sel42_b28/or_B2_B3_o ;
  wire \picorv32_core/sel42_b28/or_B4_B5_o ;
  wire \picorv32_core/sel42_b28/or_B6_B7_o ;
  wire \picorv32_core/sel42_b28/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b28/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b29/or_B0_B1_o ;
  wire \picorv32_core/sel42_b29/or_B2_B3_o ;
  wire \picorv32_core/sel42_b29/or_B4_B5_o ;
  wire \picorv32_core/sel42_b29/or_B6_B7_o ;
  wire \picorv32_core/sel42_b29/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b29/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b3/or_B0_B1_o ;
  wire \picorv32_core/sel42_b3/or_B2_B3_o ;
  wire \picorv32_core/sel42_b3/or_B4_B5_o ;
  wire \picorv32_core/sel42_b3/or_B6_B7_o ;
  wire \picorv32_core/sel42_b3/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b3/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b30/or_B0_B1_o ;
  wire \picorv32_core/sel42_b30/or_B2_B3_o ;
  wire \picorv32_core/sel42_b30/or_B4_B5_o ;
  wire \picorv32_core/sel42_b30/or_B6_B7_o ;
  wire \picorv32_core/sel42_b30/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b30/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b31/or_B0_B1_o ;
  wire \picorv32_core/sel42_b31/or_B2_B3_o ;
  wire \picorv32_core/sel42_b31/or_B4_B5_o ;
  wire \picorv32_core/sel42_b31/or_B6_B7_o ;
  wire \picorv32_core/sel42_b31/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b31/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b4/or_B0_B1_o ;
  wire \picorv32_core/sel42_b4/or_B2_B3_o ;
  wire \picorv32_core/sel42_b4/or_B4_B5_o ;
  wire \picorv32_core/sel42_b4/or_B6_B7_o ;
  wire \picorv32_core/sel42_b4/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b4/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b5/or_B0_B1_o ;
  wire \picorv32_core/sel42_b5/or_B2_B3_o ;
  wire \picorv32_core/sel42_b5/or_B4_B5_o ;
  wire \picorv32_core/sel42_b5/or_B6_B7_o ;
  wire \picorv32_core/sel42_b5/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b5/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b6/or_B0_B1_o ;
  wire \picorv32_core/sel42_b6/or_B2_B3_o ;
  wire \picorv32_core/sel42_b6/or_B4_B5_o ;
  wire \picorv32_core/sel42_b6/or_B6_B7_o ;
  wire \picorv32_core/sel42_b6/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b6/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b7/or_B0_B1_o ;
  wire \picorv32_core/sel42_b7/or_B2_B3_o ;
  wire \picorv32_core/sel42_b7/or_B4_B5_o ;
  wire \picorv32_core/sel42_b7/or_B6_B7_o ;
  wire \picorv32_core/sel42_b7/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b7/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b8/or_B0_B1_o ;
  wire \picorv32_core/sel42_b8/or_B2_B3_o ;
  wire \picorv32_core/sel42_b8/or_B4_B5_o ;
  wire \picorv32_core/sel42_b8/or_B6_B7_o ;
  wire \picorv32_core/sel42_b8/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b8/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel42_b9/or_B0_B1_o ;
  wire \picorv32_core/sel42_b9/or_B2_B3_o ;
  wire \picorv32_core/sel42_b9/or_B4_B5_o ;
  wire \picorv32_core/sel42_b9/or_B6_B7_o ;
  wire \picorv32_core/sel42_b9/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel42_b9/or_or_B4_B5_o_or_B6__o ;
  wire \picorv32_core/sel43_b0/or_B2_B3_o ;
  wire \picorv32_core/sel43_b0/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b1/or_B2_B3_o ;
  wire \picorv32_core/sel43_b1/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b10/or_B2_B3_o ;
  wire \picorv32_core/sel43_b10/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b11/or_B2_B3_o ;
  wire \picorv32_core/sel43_b11/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b12/or_B2_B3_o ;
  wire \picorv32_core/sel43_b12/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b13/or_B2_B3_o ;
  wire \picorv32_core/sel43_b13/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b14/or_B2_B3_o ;
  wire \picorv32_core/sel43_b14/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b15/or_B2_B3_o ;
  wire \picorv32_core/sel43_b15/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b16/or_B2_B3_o ;
  wire \picorv32_core/sel43_b16/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b17/or_B2_B3_o ;
  wire \picorv32_core/sel43_b17/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b18/or_B2_B3_o ;
  wire \picorv32_core/sel43_b18/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b19/or_B2_B3_o ;
  wire \picorv32_core/sel43_b19/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b2/or_B2_B3_o ;
  wire \picorv32_core/sel43_b2/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b20/or_B2_B3_o ;
  wire \picorv32_core/sel43_b20/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b21/or_B2_B3_o ;
  wire \picorv32_core/sel43_b21/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b22/or_B2_B3_o ;
  wire \picorv32_core/sel43_b22/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b23/or_B2_B3_o ;
  wire \picorv32_core/sel43_b23/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b24/or_B2_B3_o ;
  wire \picorv32_core/sel43_b24/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b25/or_B2_B3_o ;
  wire \picorv32_core/sel43_b25/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b26/or_B2_B3_o ;
  wire \picorv32_core/sel43_b26/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b27/or_B2_B3_o ;
  wire \picorv32_core/sel43_b27/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b28/or_B2_B3_o ;
  wire \picorv32_core/sel43_b28/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b29/or_B2_B3_o ;
  wire \picorv32_core/sel43_b29/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b3/or_B2_B3_o ;
  wire \picorv32_core/sel43_b3/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b30/or_B2_B3_o ;
  wire \picorv32_core/sel43_b30/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b31/or_B2_B3_o ;
  wire \picorv32_core/sel43_b31/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b4/or_B2_B3_o ;
  wire \picorv32_core/sel43_b4/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b5/or_B2_B3_o ;
  wire \picorv32_core/sel43_b5/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b6/or_B2_B3_o ;
  wire \picorv32_core/sel43_b6/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b7/or_B2_B3_o ;
  wire \picorv32_core/sel43_b7/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b8/or_B2_B3_o ;
  wire \picorv32_core/sel43_b8/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel43_b9/or_B2_B3_o ;
  wire \picorv32_core/sel43_b9/or_or_B0_B1_o_or_B2__o ;
  wire \picorv32_core/sel44_b0/or_B4_B5_o ;
  wire \picorv32_core/sel44_b1/or_B4_B5_o ;
  wire \picorv32_core/sel44_b2/or_B4_B5_o ;
  wire \picorv32_core/sel44_b3/or_B4_B5_o ;
  wire \picorv32_core/sel44_b4/or_B4_B5_o ;
  wire \picorv32_core/sel45/or_B0_B1_o ;
  wire \picorv32_core/sel45/or_B2_B3_o ;
  wire \picorv32_core/sel46_sel_is_2_o ;
  wire \picorv32_core/sel4_b0/or_B0_B1_o ;
  wire \picorv32_core/sel4_b1/or_B0_B1_o ;
  wire \picorv32_core/sel4_b2/or_B0_B1_o ;
  wire \picorv32_core/sel5_b2/or_B1_B2_o ;
  wire \picorv32_core/sel5_b3/or_B1_B2_o ;
  wire \picorv32_core/sel5_b4/or_B1_B2_o ;
  wire \picorv32_core/sel6_b1/or_B1_B2_o ;
  wire \picorv32_core/sel7/or_B1_B2_o ;
  wire \picorv32_core/u170_sel_is_2_o ;
  wire \picorv32_core/u173_sel_is_3_o ;
  wire \picorv32_core/u179_sel_is_0_o ;
  wire \picorv32_core/u235_sel_is_0_o_neg ;
  wire \picorv32_core/u239_sel_is_0_o_neg ;
  wire \picorv32_core/u247_sel_is_1_o ;
  wire \picorv32_core/u248_sel_is_1_o ;
  wire \picorv32_core/u252_sel_is_3_o ;
  wire \picorv32_core/u255_sel_is_3_o ;
  wire \picorv32_core/u256_sel_is_3_o ;
  wire \picorv32_core/u257_sel_is_3_o ;
  wire \picorv32_core/u449_sel_is_0_o ;
  wire \picorv32_core/u527_sel_is_3_o ;
  wire \picorv32_core/u589_sel_is_3_o ;
  wire \picorv32_core/u596_sel_is_3_o ;
  wire \picorv32_core/u597_sel_is_3_o ;
  wire \picorv32_core/u599_sel_is_3_o ;
  wire \picorv32_core/u616_sel_is_2_o ;
  wire \picorv32_core/u617_sel_is_2_o ;
  wire \picorv32_core/u623_sel_is_2_o ;
  wire \picorv32_core/u624_sel_is_2_o ;
  wire \picorv32_core/u625_sel_is_2_o ;
  wire \picorv32_core/u626_sel_is_2_o ;
  wire resetn;  // ../src/top.v(33)
  wire \uart/mux10_b0_sel_is_3_o ;
  wire \uart/mux12_b0_sel_is_3_o ;
  wire \uart/mux13_b0_sel_is_3_o ;
  wire \uart/mux14_b0_sel_is_1_o ;
  wire \uart/mux15_b0_sel_is_2_o ;
  wire \uart/mux37_b0_sel_is_3_o ;
  wire \uart/mux44_b0_sel_is_26_o ;
  wire \uart/mux4_sel_is_3_o ;
  wire \uart/mux51_b0_sel_is_3_o ;
  wire \uart/mux5_b0_sel_is_2_o ;
  wire \uart/mux6_b0_sel_is_4_o ;
  wire \uart/mux9_b0_sel_is_3_o ;
  wire \uart/n0 ;
  wire \uart/n112 ;
  wire \uart/n2 ;
  wire \uart/n29 ;
  wire \uart/n3 ;
  wire \uart/n30 ;
  wire \uart/n34 ;
  wire \uart/n39 ;
  wire \uart/n43 ;
  wire \uart/n44 ;
  wire \uart/n51 ;
  wire \uart/n52 ;
  wire \uart/n56 ;
  wire \uart/n58 ;
  wire \uart/n60 ;
  wire \uart/n62 ;
  wire \uart/n64 ;
  wire \uart/n66 ;
  wire \uart/n68 ;
  wire \uart/n70 ;
  wire \uart/n72 ;
  wire \uart/n74 ;
  wire \uart/n82 ;
  wire \uart/n83 ;
  wire \uart/n84 ;
  wire \uart/n85 ;
  wire \uart/n86 ;
  wire \uart/n87 ;
  wire \uart/n88 ;
  wire \uart/n89 ;
  wire \uart/n9 ;
  wire \uart/n90 ;
  wire \uart/n91 ;
  wire \uart/n96 ;
  wire \uart/n97 ;
  wire \uart/n98 ;
  wire \uart/n99 ;
  wire \uart/u7_sel_is_3_o ;
  wire \uart/u9_sel_is_3_o ;
  wire \uart/uart_op_clock ;  // ../src/uart.v(34)
  wire \uart/uart_op_clock_by_3 ;  // ../src/uart.v(37)
  wire \uart/uart_status_fe ;  // ../src/uart.v(39)
  wire \uart/uart_status_rx ;  // ../src/uart.v(40)
  wire \uart/uart_status_rx_clr ;  // ../src/uart.v(156)
  wire \uart/uart_status_rxd$0$_neg ;
  wire \uart/uart_status_rxd$2$_neg ;
  wire \uart/uart_trigger_tx ;  // ../src/uart.v(44)
  wire uart_sel;  // ../src/top.v(97)

  add_pu2_pu2_o2 add0 (
    .i0(initial_reset),
    .i1(2'b01),
    .o(n3));  // ../src/top.v(41)
  eq_w2 eq0 (
    .i0(initial_reset),
    .i1(2'b11),
    .o(n0));  // ../src/top.v(38)
  eq_w20 eq1 (
    .i0(mem_la_addr[31:12]),
    .i1(20'b00000000000000000000),
    .o(n6));  // ../src/top.v(74)
  eq_w28 eq2 (
    .i0(mem_la_addr[31:4]),
    .i1(28'b0001000000000000000000000001),
    .o(uart_sel));  // ../src/top.v(97)
  eq_w30 eq3 (
    .i0(mem_la_addr[31:2]),
    .i1(30'b000100000000000000000000000000),
    .o(n15));  // ../src/top.v(124)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("hi.mif"),
    .ADDR_WIDTH_A(10),
    .ADDR_WIDTH_B(10),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(1024),
    .DATA_DEPTH_B(1024),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .PACKABLE("NO"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \mem_hi/inst  (
    .addra(mem_la_addr[11:2]),
    .addrb(10'b0000000000),
    .bea(1'b0),
    .beb(1'b0),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(mem_la_wdata[31:24]),
    .dib(8'b00000000),
    .ocea(1'b0),
    .oceb(1'b0),
    .rsta(\picorv32_core/n407 ),
    .rstb(1'b0),
    .wea(n13),
    .web(1'b0),
    .doa(memory_out[31:24]));  // al_ip/mem_hi.v(43)
  not \mem_la_addr[2]_inv  (mem_la_addr$2$_neg, mem_la_addr[2]);
  not \mem_la_addr[3]_inv  (mem_la_addr$3$_neg, mem_la_addr[3]);
  not mem_la_write_inv (mem_la_write_neg, mem_la_write);
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("lo.mif"),
    .ADDR_WIDTH_A(10),
    .ADDR_WIDTH_B(10),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(1024),
    .DATA_DEPTH_B(1024),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .PACKABLE("NO"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \mem_lo/inst  (
    .addra(mem_la_addr[11:2]),
    .addrb(10'b0000000000),
    .bea(1'b0),
    .beb(1'b0),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(mem_la_wdata[7:0]),
    .dib(8'b00000000),
    .ocea(1'b0),
    .oceb(1'b0),
    .rsta(\picorv32_core/n407 ),
    .rstb(1'b0),
    .wea(n7),
    .web(1'b0),
    .doa(memory_out[7:0]));  // al_ip/mem_lo.v(43)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("mh.mif"),
    .ADDR_WIDTH_A(10),
    .ADDR_WIDTH_B(10),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(1024),
    .DATA_DEPTH_B(1024),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .PACKABLE("NO"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \mem_mh/inst  (
    .addra(mem_la_addr[11:2]),
    .addrb(10'b0000000000),
    .bea(1'b0),
    .beb(1'b0),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(mem_la_wdata[23:16]),
    .dib(8'b00000000),
    .ocea(1'b0),
    .oceb(1'b0),
    .rsta(\picorv32_core/n407 ),
    .rstb(1'b0),
    .wea(n11),
    .web(1'b0),
    .doa(memory_out[23:16]));  // al_ip/mem_mh.v(43)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("ml.mif"),
    .ADDR_WIDTH_A(10),
    .ADDR_WIDTH_B(10),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(1024),
    .DATA_DEPTH_B(1024),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .PACKABLE("NO"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \mem_ml/inst  (
    .addra(mem_la_addr[11:2]),
    .addrb(10'b0000000000),
    .bea(1'b0),
    .beb(1'b0),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(mem_la_wdata[15:8]),
    .dib(8'b00000000),
    .ocea(1'b0),
    .oceb(1'b0),
    .rsta(\picorv32_core/n407 ),
    .rstb(1'b0),
    .wea(n9),
    .web(1'b0),
    .doa(memory_out[15:8]));  // al_ip/mem_ml.v(43)
  binary_mux_s1_w1 mux1_b0 (
    .i0(memory_out[0]),
    .i1(uart_do[0]),
    .sel(uart_sel),
    .o(mem_rdata[0]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b1 (
    .i0(memory_out[1]),
    .i1(uart_do[1]),
    .sel(uart_sel),
    .o(mem_rdata[1]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b10 (
    .i0(memory_out[10]),
    .i1(uart_do[10]),
    .sel(uart_sel),
    .o(mem_rdata[10]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b11 (
    .i0(memory_out[11]),
    .i1(uart_do[11]),
    .sel(uart_sel),
    .o(mem_rdata[11]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b12 (
    .i0(memory_out[12]),
    .i1(uart_do[12]),
    .sel(uart_sel),
    .o(mem_rdata[12]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b13 (
    .i0(memory_out[13]),
    .i1(uart_do[13]),
    .sel(uart_sel),
    .o(mem_rdata[13]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b14 (
    .i0(memory_out[14]),
    .i1(uart_do[14]),
    .sel(uart_sel),
    .o(mem_rdata[14]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b15 (
    .i0(memory_out[15]),
    .i1(uart_do[15]),
    .sel(uart_sel),
    .o(mem_rdata[15]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b16 (
    .i0(memory_out[16]),
    .i1(uart_do[16]),
    .sel(uart_sel),
    .o(mem_rdata[16]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b17 (
    .i0(memory_out[17]),
    .i1(uart_do[17]),
    .sel(uart_sel),
    .o(mem_rdata[17]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b18 (
    .i0(memory_out[18]),
    .i1(uart_do[18]),
    .sel(uart_sel),
    .o(mem_rdata[18]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b19 (
    .i0(memory_out[19]),
    .i1(uart_do[19]),
    .sel(uart_sel),
    .o(mem_rdata[19]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b2 (
    .i0(memory_out[2]),
    .i1(uart_do[2]),
    .sel(uart_sel),
    .o(mem_rdata[2]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b20 (
    .i0(memory_out[20]),
    .i1(uart_do[20]),
    .sel(uart_sel),
    .o(mem_rdata[20]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b21 (
    .i0(memory_out[21]),
    .i1(uart_do[21]),
    .sel(uart_sel),
    .o(mem_rdata[21]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b22 (
    .i0(memory_out[22]),
    .i1(uart_do[22]),
    .sel(uart_sel),
    .o(mem_rdata[22]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b23 (
    .i0(memory_out[23]),
    .i1(uart_do[23]),
    .sel(uart_sel),
    .o(mem_rdata[23]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b24 (
    .i0(memory_out[24]),
    .i1(uart_do[24]),
    .sel(uart_sel),
    .o(mem_rdata[24]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b25 (
    .i0(memory_out[25]),
    .i1(uart_do[25]),
    .sel(uart_sel),
    .o(mem_rdata[25]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b26 (
    .i0(memory_out[26]),
    .i1(uart_do[26]),
    .sel(uart_sel),
    .o(mem_rdata[26]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b27 (
    .i0(memory_out[27]),
    .i1(uart_do[27]),
    .sel(uart_sel),
    .o(mem_rdata[27]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b28 (
    .i0(memory_out[28]),
    .i1(uart_do[28]),
    .sel(uart_sel),
    .o(mem_rdata[28]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b29 (
    .i0(memory_out[29]),
    .i1(uart_do[29]),
    .sel(uart_sel),
    .o(mem_rdata[29]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b3 (
    .i0(memory_out[3]),
    .i1(uart_do[3]),
    .sel(uart_sel),
    .o(mem_rdata[3]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b30 (
    .i0(memory_out[30]),
    .i1(uart_do[30]),
    .sel(uart_sel),
    .o(mem_rdata[30]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b31 (
    .i0(memory_out[31]),
    .i1(uart_do[31]),
    .sel(uart_sel),
    .o(mem_rdata[31]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b4 (
    .i0(memory_out[4]),
    .i1(uart_do[4]),
    .sel(uart_sel),
    .o(mem_rdata[4]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b5 (
    .i0(memory_out[5]),
    .i1(uart_do[5]),
    .sel(uart_sel),
    .o(mem_rdata[5]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b6 (
    .i0(memory_out[6]),
    .i1(uart_do[6]),
    .sel(uart_sel),
    .o(mem_rdata[6]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b7 (
    .i0(memory_out[7]),
    .i1(uart_do[7]),
    .sel(uart_sel),
    .o(mem_rdata[7]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b8 (
    .i0(memory_out[8]),
    .i1(uart_do[8]),
    .sel(uart_sel),
    .o(mem_rdata[8]));  // ../src/top.v(110)
  binary_mux_s1_w1 mux1_b9 (
    .i0(memory_out[9]),
    .i1(uart_do[9]),
    .sel(uart_sel),
    .o(mem_rdata[9]));  // ../src/top.v(110)
  ne_w2 neq0 (
    .i0(initial_reset),
    .i1(2'b11),
    .o(n2));  // ../src/top.v(40)
  reg_ar_as_w1 out_byte_en_reg (
    .clk(clk),
    .d(n16),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(out_byte_en));  // ../src/top.v(128)
  add_pu30_pu30_o30 \picorv32_core/add0  (
    .i0(\picorv32_core/next_pc [31:2]),
    .i1({29'b00000000000000000000000000000,\picorv32_core/mem_la_firstword_xfer }),
    .o(\picorv32_core/n30 ));  // ../src/picorv32.v(346)
  add_pu32_pu32_o32 \picorv32_core/add1  (
    .i0({\picorv32_core/pcpi_rs1$31$ ,\picorv32_core/pcpi_rs1$30$ ,\picorv32_core/pcpi_rs1$29$ ,\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$25$ ,\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/pcpi_rs1$23$ ,\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs1$21$ ,\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/pcpi_rs1$19$ ,\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$17$ ,\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/pcpi_rs1$15$ ,\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/pcpi_rs1$11$ ,\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$9$ ,\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/pcpi_rs1$7$ ,\picorv32_core/pcpi_rs1$6$ ,\picorv32_core/pcpi_rs1$5$ ,\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/pcpi_rs1$3$ ,\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .i1({\picorv32_core/pcpi_rs2$31$ ,\picorv32_core/pcpi_rs2$30$ ,\picorv32_core/pcpi_rs2$29$ ,\picorv32_core/pcpi_rs2$28$ ,\picorv32_core/pcpi_rs2$27$ ,\picorv32_core/pcpi_rs2$26$ ,\picorv32_core/pcpi_rs2$25$ ,\picorv32_core/pcpi_rs2$24$ ,\picorv32_core/pcpi_rs2$23$ ,\picorv32_core/pcpi_rs2$22$ ,\picorv32_core/pcpi_rs2$21$ ,\picorv32_core/pcpi_rs2$20$ ,\picorv32_core/pcpi_rs2$19$ ,\picorv32_core/pcpi_rs2$18$ ,\picorv32_core/pcpi_rs2$17$ ,\picorv32_core/pcpi_rs2$16$ ,\picorv32_core/pcpi_rs2$15$ ,\picorv32_core/pcpi_rs2$14$ ,\picorv32_core/pcpi_rs2$13$ ,\picorv32_core/pcpi_rs2$12$ ,\picorv32_core/pcpi_rs2$11$ ,\picorv32_core/pcpi_rs2$10$ ,\picorv32_core/pcpi_rs2$9$ ,\picorv32_core/pcpi_rs2$8$ ,mem_la_wdata[7:0]}),
    .o(\picorv32_core/n434 ));  // ../src/picorv32.v(1193)
  add_pu32_pu32_o32 \picorv32_core/add2  (
    .i0(\picorv32_core/reg_pc ),
    .i1({29'b00000000000000000000000000000,\picorv32_core/n449 [2],\picorv32_core/latched_compr ,1'b0}),
    .o(\picorv32_core/n450 ));  // ../src/picorv32.v(1270)
  add_pu64_pu64_o64 \picorv32_core/add3  (
    .i0(\picorv32_core/count_cycle ),
    .i1(64'b0000000000000000000000000000000000000000000000000000000000000001),
    .o(\picorv32_core/n459 ));  // ../src/picorv32.v(1365)
  add_pu32_pu32_o32 \picorv32_core/add4  (
    .i0(\picorv32_core/n500 ),
    .i1({29'b00000000000000000000000000000,\picorv32_core/n501 [2],\picorv32_core/compressed_instr ,1'b0}),
    .o(\picorv32_core/n502 ));  // ../src/picorv32.v(1498)
  add_pu64_pu64_o64 \picorv32_core/add5  (
    .i0(\picorv32_core/count_instr ),
    .i1(64'b0000000000000000000000000000000000000000000000000000000000000001),
    .o(\picorv32_core/n503 ));  // ../src/picorv32.v(1502)
  add_pu32_pu32_o32 \picorv32_core/add6  (
    .i0(\picorv32_core/n500 ),
    .i1({\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20],\picorv32_core/decoded_imm_uj [20:1],1'b0}),
    .o(\picorv32_core/n504 ));  // ../src/picorv32.v(1507)
  add_pu32_pu32_o32 \picorv32_core/add7  (
    .i0(\picorv32_core/reg_pc ),
    .i1(\picorv32_core/decoded_imm ),
    .o(\picorv32_core/n543 ));  // ../src/picorv32.v(1744)
  add_pu32_pu32_o32 \picorv32_core/add8  (
    .i0({\picorv32_core/pcpi_rs1$31$ ,\picorv32_core/pcpi_rs1$30$ ,\picorv32_core/pcpi_rs1$29$ ,\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$25$ ,\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/pcpi_rs1$23$ ,\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs1$21$ ,\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/pcpi_rs1$19$ ,\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$17$ ,\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/pcpi_rs1$15$ ,\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/pcpi_rs1$11$ ,\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$9$ ,\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/pcpi_rs1$7$ ,\picorv32_core/pcpi_rs1$6$ ,\picorv32_core/pcpi_rs1$5$ ,\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/pcpi_rs1$3$ ,\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .i1(\picorv32_core/decoded_imm ),
    .o(\picorv32_core/n576 ));  // ../src/picorv32.v(1807)
  not \picorv32_core/clear_prefetched_high_word_inv  (\picorv32_core/clear_prefetched_high_word_neg , \picorv32_core/clear_prefetched_high_word );
  reg_ar_ss_w1 \picorv32_core/clear_prefetched_high_word_q_reg  (
    .clk(clk),
    .d(1'b0),
    .en(~\picorv32_core/prefetched_high_word ),
    .reset(1'b0),
    .set(\picorv32_core/n447 ),
    .q(\picorv32_core/clear_prefetched_high_word_q ));  // ../src/picorv32.v(1241)
  reg_ar_as_w1 \picorv32_core/compressed_instr_reg  (
    .clk(clk),
    .d(\picorv32_core/n180 ),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/compressed_instr ));  // ../src/picorv32.v(1120)
  EG_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(32),
    .DATA_WIDTH_W(32),
    .INIT_FILE("zero.mif"))
    \picorv32_core/cpuregs_p1/dram  (
    .di(\picorv32_core/cpuregs_wrdata ),
    .raddr(\picorv32_core/decoded_rs1 ),
    .waddr(\picorv32_core/latched_rd ),
    .wclk(clk),
    .we(\picorv32_core/n456 ),
    .do(\picorv32_core/cpuregs_rs1_z ));  // al_ip/cpuregs.v(40)
  EG_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(32),
    .DATA_WIDTH_W(32),
    .INIT_FILE("zero.mif"))
    \picorv32_core/cpuregs_p2/dram  (
    .di(\picorv32_core/cpuregs_wrdata ),
    .raddr(\picorv32_core/decoded_rs2 ),
    .waddr(\picorv32_core/latched_rd ),
    .wclk(clk),
    .we(\picorv32_core/n456 ),
    .do(\picorv32_core/cpuregs_rs2_z ));  // al_ip/cpuregs.v(40)
  reg_sr_as_w1 \picorv32_core/decoder_pseudo_trigger_reg  (
    .clk(clk),
    .d(\picorv32_core/n580 ),
    .en(1'b1),
    .reset(~\picorv32_core/u625_sel_is_2_o ),
    .set(1'b0),
    .q(\picorv32_core/decoder_pseudo_trigger ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/decoder_trigger_reg  (
    .clk(clk),
    .d(\picorv32_core/n727 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoder_trigger ));  // ../src/picorv32.v(1906)
  eq_w3 \picorv32_core/eq0  (
    .i0(\picorv32_core/mem_rdata_latched [15:13]),
    .i1(3'b000),
    .o(\picorv32_core/n96 ));  // ../src/picorv32.v(404)
  eq_w3 \picorv32_core/eq1  (
    .i0(\picorv32_core/mem_rdata_latched [15:13]),
    .i1(3'b010),
    .o(\picorv32_core/n97 ));  // ../src/picorv32.v(408)
  eq_w2 \picorv32_core/eq10  (
    .i0(\picorv32_core/mem_rdata_latched [6:5]),
    .i1(2'b10),
    .o(\picorv32_core/n65 ));  // ../src/picorv32.v(453)
  eq_w2 \picorv32_core/eq11  (
    .i0(\picorv32_core/mem_rdata_latched [6:5]),
    .i1(2'b11),
    .o(\picorv32_core/n67 ));  // ../src/picorv32.v(454)
  eq_w1 \picorv32_core/eq12  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(1'b0),
    .o(\picorv32_core/n72 ));  // ../src/picorv32.v(483)
  eq_w5 \picorv32_core/eq13  (
    .i0(\picorv32_core/mem_rdata_latched [6:2]),
    .i1(5'b00000),
    .o(\picorv32_core/n73 ));  // ../src/picorv32.v(483)
  eq_w3 \picorv32_core/eq14  (
    .i0(\picorv32_core/mem_rdata_latched [15:13]),
    .i1(3'b100),
    .o(\picorv32_core/n98 ));  // ../src/picorv32.v(482)
  eq_w7 \picorv32_core/eq15  (
    .i0(\picorv32_core/mem_rdata_latched [6:0]),
    .i1(7'b0110111),
    .o(\picorv32_core/n171 ));  // ../src/picorv32.v(829)
  eq_w7 \picorv32_core/eq16  (
    .i0(\picorv32_core/mem_rdata_latched [6:0]),
    .i1(7'b0010111),
    .o(\picorv32_core/n172 ));  // ../src/picorv32.v(830)
  eq_w7 \picorv32_core/eq17  (
    .i0(\picorv32_core/mem_rdata_latched [6:0]),
    .i1(7'b1101111),
    .o(\picorv32_core/n173 ));  // ../src/picorv32.v(831)
  eq_w7 \picorv32_core/eq18  (
    .i0(\picorv32_core/mem_rdata_latched [6:0]),
    .i1(7'b1100111),
    .o(\picorv32_core/n174 ));  // ../src/picorv32.v(832)
  eq_w7 \picorv32_core/eq19  (
    .i0(\picorv32_core/mem_rdata_latched [6:0]),
    .i1(7'b1100011),
    .o(\picorv32_core/n175 ));  // ../src/picorv32.v(836)
  eq_w3 \picorv32_core/eq2  (
    .i0(\picorv32_core/mem_rdata_latched [15:13]),
    .i1(3'b110),
    .o(\picorv32_core/n99 ));  // ../src/picorv32.v(412)
  eq_w7 \picorv32_core/eq20  (
    .i0(\picorv32_core/mem_rdata_latched [6:0]),
    .i1(7'b0000011),
    .o(\picorv32_core/n176 ));  // ../src/picorv32.v(837)
  eq_w7 \picorv32_core/eq21  (
    .i0(\picorv32_core/mem_rdata_latched [6:0]),
    .i1(7'b0100011),
    .o(\picorv32_core/n177 ));  // ../src/picorv32.v(838)
  eq_w7 \picorv32_core/eq22  (
    .i0(\picorv32_core/mem_rdata_latched [6:0]),
    .i1(7'b0010011),
    .o(\picorv32_core/n178 ));  // ../src/picorv32.v(839)
  eq_w7 \picorv32_core/eq23  (
    .i0(\picorv32_core/mem_rdata_latched [6:0]),
    .i1(7'b0110011),
    .o(\picorv32_core/n179 ));  // ../src/picorv32.v(840)
  eq_w3 \picorv32_core/eq24  (
    .i0(\picorv32_core/mem_rdata_q [14:12]),
    .i1(3'b000),
    .o(\picorv32_core/n275 ));  // ../src/picorv32.v(996)
  eq_w3 \picorv32_core/eq25  (
    .i0(\picorv32_core/mem_rdata_q [14:12]),
    .i1(3'b001),
    .o(\picorv32_core/n277 ));  // ../src/picorv32.v(997)
  eq_w3 \picorv32_core/eq26  (
    .i0(\picorv32_core/mem_rdata_q [14:12]),
    .i1(3'b100),
    .o(\picorv32_core/n279 ));  // ../src/picorv32.v(998)
  eq_w3 \picorv32_core/eq27  (
    .i0(\picorv32_core/mem_rdata_q [14:12]),
    .i1(3'b101),
    .o(\picorv32_core/n281 ));  // ../src/picorv32.v(999)
  eq_w3 \picorv32_core/eq28  (
    .i0(\picorv32_core/mem_rdata_q [14:12]),
    .i1(3'b110),
    .o(\picorv32_core/n283 ));  // ../src/picorv32.v(1000)
  eq_w3 \picorv32_core/eq29  (
    .i0(\picorv32_core/mem_rdata_q [14:12]),
    .i1(3'b111),
    .o(\picorv32_core/n285 ));  // ../src/picorv32.v(1001)
  eq_w5 \picorv32_core/eq3  (
    .i0(\picorv32_core/mem_rdata_latched [11:7]),
    .i1(5'b00010),
    .o(\picorv32_core/n193 ));  // ../src/picorv32.v(429)
  eq_w3 \picorv32_core/eq30  (
    .i0(\picorv32_core/mem_rdata_q [14:12]),
    .i1(3'b010),
    .o(\picorv32_core/n289 ));  // ../src/picorv32.v(1005)
  eq_w3 \picorv32_core/eq31  (
    .i0(\picorv32_core/mem_rdata_q [14:12]),
    .i1(3'b011),
    .o(\picorv32_core/n298 ));  // ../src/picorv32.v(1015)
  eq_w7 \picorv32_core/eq32  (
    .i0(\picorv32_core/mem_rdata_q [31:25]),
    .i1(7'b0000000),
    .o(\picorv32_core/n304 ));  // ../src/picorv32.v(1020)
  eq_w7 \picorv32_core/eq33  (
    .i0(\picorv32_core/mem_rdata_q [31:25]),
    .i1(7'b0100000),
    .o(\picorv32_core/n308 ));  // ../src/picorv32.v(1022)
  eq_w7 \picorv32_core/eq34  (
    .i0(\picorv32_core/mem_rdata_q [6:0]),
    .i1(7'b1110011),
    .o(\picorv32_core/n328 ));  // ../src/picorv32.v(1035)
  eq_w20 \picorv32_core/eq35  (
    .i0(\picorv32_core/mem_rdata_q [31:12]),
    .i1(20'b11000000000000000010),
    .o(\picorv32_core/n329 ));  // ../src/picorv32.v(1035)
  eq_w20 \picorv32_core/eq36  (
    .i0(\picorv32_core/mem_rdata_q [31:12]),
    .i1(20'b11000000000100000010),
    .o(\picorv32_core/n331 ));  // ../src/picorv32.v(1036)
  eq_w20 \picorv32_core/eq37  (
    .i0(\picorv32_core/mem_rdata_q [31:12]),
    .i1(20'b11001000000000000010),
    .o(\picorv32_core/n334 ));  // ../src/picorv32.v(1037)
  eq_w20 \picorv32_core/eq38  (
    .i0(\picorv32_core/mem_rdata_q [31:12]),
    .i1(20'b11001000000100000010),
    .o(\picorv32_core/n336 ));  // ../src/picorv32.v(1038)
  eq_w20 \picorv32_core/eq39  (
    .i0(\picorv32_core/mem_rdata_q [31:12]),
    .i1(20'b11000000001000000010),
    .o(\picorv32_core/n339 ));  // ../src/picorv32.v(1039)
  eq_w2 \picorv32_core/eq4  (
    .i0(\picorv32_core/mem_rdata_latched [11:10]),
    .i1(2'b00),
    .o(\picorv32_core/n54 ));  // ../src/picorv32.v(438)
  eq_w20 \picorv32_core/eq40  (
    .i0(\picorv32_core/mem_rdata_q [31:12]),
    .i1(20'b11001000001000000010),
    .o(\picorv32_core/n341 ));  // ../src/picorv32.v(1040)
  eq_w32 \picorv32_core/eq41  (
    .i0({\picorv32_core/pcpi_rs1$31$ ,\picorv32_core/pcpi_rs1$30$ ,\picorv32_core/pcpi_rs1$29$ ,\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$25$ ,\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/pcpi_rs1$23$ ,\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs1$21$ ,\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/pcpi_rs1$19$ ,\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$17$ ,\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/pcpi_rs1$15$ ,\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/pcpi_rs1$11$ ,\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$9$ ,\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/pcpi_rs1$7$ ,\picorv32_core/pcpi_rs1$6$ ,\picorv32_core/pcpi_rs1$5$ ,\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/pcpi_rs1$3$ ,\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .i1({\picorv32_core/pcpi_rs2$31$ ,\picorv32_core/pcpi_rs2$30$ ,\picorv32_core/pcpi_rs2$29$ ,\picorv32_core/pcpi_rs2$28$ ,\picorv32_core/pcpi_rs2$27$ ,\picorv32_core/pcpi_rs2$26$ ,\picorv32_core/pcpi_rs2$25$ ,\picorv32_core/pcpi_rs2$24$ ,\picorv32_core/pcpi_rs2$23$ ,\picorv32_core/pcpi_rs2$22$ ,\picorv32_core/pcpi_rs2$21$ ,\picorv32_core/pcpi_rs2$20$ ,\picorv32_core/pcpi_rs2$19$ ,\picorv32_core/pcpi_rs2$18$ ,\picorv32_core/pcpi_rs2$17$ ,\picorv32_core/pcpi_rs2$16$ ,\picorv32_core/pcpi_rs2$15$ ,\picorv32_core/pcpi_rs2$14$ ,\picorv32_core/pcpi_rs2$13$ ,\picorv32_core/pcpi_rs2$12$ ,\picorv32_core/pcpi_rs2$11$ ,\picorv32_core/pcpi_rs2$10$ ,\picorv32_core/pcpi_rs2$9$ ,\picorv32_core/pcpi_rs2$8$ ,mem_la_wdata[7:0]}),
    .o(\picorv32_core/alu_eq ));  // ../src/picorv32.v(1194)
  eq_w8 \picorv32_core/eq42  (
    .i0(\picorv32_core/cpu_state ),
    .i1(8'b01000000),
    .o(\picorv32_core/n663 ));  // ../src/picorv32.v(1266)
  eq_w5 \picorv32_core/eq43  (
    .i0(\picorv32_core/reg_sh ),
    .i1(5'b00000),
    .o(\picorv32_core/n553 ));  // ../src/picorv32.v(1769)
  eq_w8 \picorv32_core/eq44  (
    .i0(\picorv32_core/cpu_state ),
    .i1(8'b10000000),
    .o(\picorv32_core/n662 ));  // ../src/picorv32.v(1425)
  eq_w8 \picorv32_core/eq45  (
    .i0(\picorv32_core/cpu_state ),
    .i1(8'b00100000),
    .o(\picorv32_core/n664 ));  // ../src/picorv32.v(1517)
  eq_w8 \picorv32_core/eq46  (
    .i0(\picorv32_core/cpu_state ),
    .i1(8'b00010000),
    .o(\picorv32_core/n665 ));  // ../src/picorv32.v(1697)
  eq_w8 \picorv32_core/eq47  (
    .i0(\picorv32_core/cpu_state ),
    .i1(8'b00001000),
    .o(\picorv32_core/n666 ));  // ../src/picorv32.v(1743)
  eq_w8 \picorv32_core/eq48  (
    .i0(\picorv32_core/cpu_state ),
    .i1(8'b00000100),
    .o(\picorv32_core/n667 ));  // ../src/picorv32.v(1767)
  eq_w8 \picorv32_core/eq49  (
    .i0(\picorv32_core/cpu_state ),
    .i1(8'b00000010),
    .o(\picorv32_core/n668 ));  // ../src/picorv32.v(1792)
  eq_w2 \picorv32_core/eq5  (
    .i0(\picorv32_core/mem_rdata_latched [11:10]),
    .i1(2'b01),
    .o(\picorv32_core/n56 ));  // ../src/picorv32.v(442)
  eq_w8 \picorv32_core/eq50  (
    .i0(\picorv32_core/cpu_state ),
    .i1(8'b00000001),
    .o(\picorv32_core/n669 ));  // ../src/picorv32.v(1818)
  eq_w2 \picorv32_core/eq51  (
    .i0(\picorv32_core/mem_wordsize ),
    .i1(2'b00),
    .o(\picorv32_core/n734 ));  // ../src/picorv32.v(1854)
  eq_w2 \picorv32_core/eq52  (
    .i0(\picorv32_core/mem_wordsize ),
    .i1(2'b01),
    .o(\picorv32_core/n738 ));  // ../src/picorv32.v(1861)
  eq_w2 \picorv32_core/eq6  (
    .i0(\picorv32_core/mem_rdata_latched [11:10]),
    .i1(2'b10),
    .o(\picorv32_core/n58 ));  // ../src/picorv32.v(446)
  eq_w3 \picorv32_core/eq7  (
    .i0(\picorv32_core/mem_rdata_latched [12:10]),
    .i1(3'b011),
    .o(\picorv32_core/n203 ));  // ../src/picorv32.v(450)
  eq_w2 \picorv32_core/eq8  (
    .i0(\picorv32_core/mem_rdata_latched [6:5]),
    .i1(2'b00),
    .o(\picorv32_core/n61 ));  // ../src/picorv32.v(451)
  eq_w2 \picorv32_core/eq9  (
    .i0(\picorv32_core/mem_rdata_latched [6:5]),
    .i1(2'b01),
    .o(\picorv32_core/n63 ));  // ../src/picorv32.v(452)
  reg_sr_as_w1 \picorv32_core/instr_add_reg  (
    .clk(clk),
    .d(\picorv32_core/n311 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_add ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_addi_reg  (
    .clk(clk),
    .d(\picorv32_core/n296 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_addi ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_and_reg  (
    .clk(clk),
    .d(\picorv32_core/n327 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_and ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_andi_reg  (
    .clk(clk),
    .d(\picorv32_core/n302 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_andi ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_auipc_reg  (
    .clk(clk),
    .d(\picorv32_core/n172 ),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_auipc ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_beq_reg  (
    .clk(clk),
    .d(\picorv32_core/n276 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_beq ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_bge_reg  (
    .clk(clk),
    .d(\picorv32_core/n282 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_bge ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_bgeu_reg  (
    .clk(clk),
    .d(\picorv32_core/n286 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_bgeu ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_blt_reg  (
    .clk(clk),
    .d(\picorv32_core/n280 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_blt ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_bltu_reg  (
    .clk(clk),
    .d(\picorv32_core/n284 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_bltu ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_bne_reg  (
    .clk(clk),
    .d(\picorv32_core/n278 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_bne ));  // ../src/picorv32.v(1120)
  not \picorv32_core/instr_jal_inv  (\picorv32_core/instr_jal_neg , \picorv32_core/instr_jal );
  reg_ar_as_w1 \picorv32_core/instr_jal_reg  (
    .clk(clk),
    .d(\picorv32_core/n255 ),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_jal ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_jalr_reg  (
    .clk(clk),
    .d(\picorv32_core/n251 ),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_jalr ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_lb_reg  (
    .clk(clk),
    .d(\picorv32_core/n287 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_lb ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_lbu_reg  (
    .clk(clk),
    .d(\picorv32_core/n291 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_lbu ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_lh_reg  (
    .clk(clk),
    .d(\picorv32_core/n288 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_lh ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_lhu_reg  (
    .clk(clk),
    .d(\picorv32_core/n292 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_lhu ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_lui_reg  (
    .clk(clk),
    .d(\picorv32_core/n256 ),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_lui ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_lw_reg  (
    .clk(clk),
    .d(\picorv32_core/n290 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_lw ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_or_reg  (
    .clk(clk),
    .d(\picorv32_core/n325 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_or ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_ori_reg  (
    .clk(clk),
    .d(\picorv32_core/n301 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_ori ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_rdcycle_reg  (
    .clk(clk),
    .d(\picorv32_core/n333 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_rdcycle ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_rdcycleh_reg  (
    .clk(clk),
    .d(\picorv32_core/n338 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_rdcycleh ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_rdinstr_reg  (
    .clk(clk),
    .d(\picorv32_core/n340 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_rdinstr ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_rdinstrh_reg  (
    .clk(clk),
    .d(\picorv32_core/n342 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_rdinstrh ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_sb_reg  (
    .clk(clk),
    .d(\picorv32_core/n293 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_sb ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_sh_reg  (
    .clk(clk),
    .d(\picorv32_core/n294 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_sh ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_sll_reg  (
    .clk(clk),
    .d(\picorv32_core/n314 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_sll ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_slli_reg  (
    .clk(clk),
    .d(\picorv32_core/n305 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_slli ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_slt_reg  (
    .clk(clk),
    .d(\picorv32_core/n316 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_slt ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_slti_reg  (
    .clk(clk),
    .d(\picorv32_core/n297 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_slti ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_sltiu_reg  (
    .clk(clk),
    .d(\picorv32_core/n299 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_sltiu ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_sltu_reg  (
    .clk(clk),
    .d(\picorv32_core/n318 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_sltu ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_sra_reg  (
    .clk(clk),
    .d(\picorv32_core/n323 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_sra ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_srai_reg  (
    .clk(clk),
    .d(\picorv32_core/n309 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_srai ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_srl_reg  (
    .clk(clk),
    .d(\picorv32_core/n322 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_srl ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_srli_reg  (
    .clk(clk),
    .d(\picorv32_core/n307 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_srli ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_sub_reg  (
    .clk(clk),
    .d(\picorv32_core/n312 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_sub ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/instr_sw_reg  (
    .clk(clk),
    .d(\picorv32_core/n295 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/instr_sw ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_xor_reg  (
    .clk(clk),
    .d(\picorv32_core/n320 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_xor ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/instr_xori_reg  (
    .clk(clk),
    .d(\picorv32_core/n300 ),
    .en(\picorv32_core/n274 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/instr_xori ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/is_alu_reg_imm_reg  (
    .clk(clk),
    .d(\picorv32_core/n249 ),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/is_alu_reg_imm ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/is_alu_reg_reg_reg  (
    .clk(clk),
    .d(\picorv32_core/n252 ),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/is_alu_reg_reg ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu_reg  (
    .clk(clk),
    .d(\picorv32_core/n254 ),
    .en(\picorv32_core/n170 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/is_compare_reg  (
    .clk(clk),
    .d(\picorv32_core/n169 ),
    .en(1'b1),
    .reset(~\picorv32_core/u449_sel_is_0_o ),
    .set(1'b0),
    .q(\picorv32_core/is_compare ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/is_jalr_addi_slti_sltiu_xori_ori_andi_reg  (
    .clk(clk),
    .d(\picorv32_core/n350 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/is_jalr_addi_slti_sltiu_xori_ori_andi ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/is_lb_lh_lw_lbu_lhu_reg  (
    .clk(clk),
    .d(\picorv32_core/n250 ),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/is_lb_lh_lw_lbu_lhu ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/is_lbu_lhu_lw_reg  (
    .clk(clk),
    .d(\picorv32_core/n168 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/is_lbu_lhu_lw ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub_reg  (
    .clk(clk),
    .d(\picorv32_core/n165 ),
    .en(1'b1),
    .reset(\picorv32_core/n274 ),
    .set(1'b0),
    .q(\picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/is_lui_auipc_jal_reg  (
    .clk(clk),
    .d(\picorv32_core/n472 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/is_lui_auipc_jal ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/is_sb_sh_sw_reg  (
    .clk(clk),
    .d(\picorv32_core/n253 ),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/is_sb_sh_sw ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/is_sll_srl_sra_reg  (
    .clk(clk),
    .d(\picorv32_core/n354 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/is_sll_srl_sra ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/is_slli_srli_srai_reg  (
    .clk(clk),
    .d(\picorv32_core/n347 ),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/is_slli_srli_srai ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/is_slti_blt_slt_reg  (
    .clk(clk),
    .d(\picorv32_core/n166 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/is_slti_blt_slt ));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/is_sltiu_bltu_sltu_reg  (
    .clk(clk),
    .d(\picorv32_core/n167 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/is_sltiu_bltu_sltu ));  // ../src/picorv32.v(1120)
  reg_sr_as_w1 \picorv32_core/latched_branch_reg  (
    .clk(clk),
    .d(\picorv32_core/n681 ),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/latched_branch ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/latched_compr_reg  (
    .clk(clk),
    .d(\picorv32_core/compressed_instr ),
    .en(\picorv32_core/u616_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/latched_compr ));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/latched_is_lb_reg  (
    .clk(clk),
    .d(\picorv32_core/n687 ),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/latched_is_lb ));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/latched_is_lh_reg  (
    .clk(clk),
    .d(\picorv32_core/n685 ),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/latched_is_lh ));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/latched_is_lu_reg  (
    .clk(clk),
    .d(\picorv32_core/n683 ),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/latched_is_lu ));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/latched_stalu_reg  (
    .clk(clk),
    .d(\picorv32_core/n679 ),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/latched_stalu ));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/latched_store_reg  (
    .clk(clk),
    .d(\picorv32_core/n677 ),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/latched_store ));  // ../src/picorv32.v(1906)
  lt_u32_u32 \picorv32_core/lt0  (
    .ci(1'b0),
    .i0({\picorv32_core/pcpi_rs2$31$ ,\picorv32_core/pcpi_rs1$30$ ,\picorv32_core/pcpi_rs1$29$ ,\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$25$ ,\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/pcpi_rs1$23$ ,\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs1$21$ ,\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/pcpi_rs1$19$ ,\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$17$ ,\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/pcpi_rs1$15$ ,\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/pcpi_rs1$11$ ,\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$9$ ,\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/pcpi_rs1$7$ ,\picorv32_core/pcpi_rs1$6$ ,\picorv32_core/pcpi_rs1$5$ ,\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/pcpi_rs1$3$ ,\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .i1({\picorv32_core/pcpi_rs1$31$ ,\picorv32_core/pcpi_rs2$30$ ,\picorv32_core/pcpi_rs2$29$ ,\picorv32_core/pcpi_rs2$28$ ,\picorv32_core/pcpi_rs2$27$ ,\picorv32_core/pcpi_rs2$26$ ,\picorv32_core/pcpi_rs2$25$ ,\picorv32_core/pcpi_rs2$24$ ,\picorv32_core/pcpi_rs2$23$ ,\picorv32_core/pcpi_rs2$22$ ,\picorv32_core/pcpi_rs2$21$ ,\picorv32_core/pcpi_rs2$20$ ,\picorv32_core/pcpi_rs2$19$ ,\picorv32_core/pcpi_rs2$18$ ,\picorv32_core/pcpi_rs2$17$ ,\picorv32_core/pcpi_rs2$16$ ,\picorv32_core/pcpi_rs2$15$ ,\picorv32_core/pcpi_rs2$14$ ,\picorv32_core/pcpi_rs2$13$ ,\picorv32_core/pcpi_rs2$12$ ,\picorv32_core/pcpi_rs2$11$ ,\picorv32_core/pcpi_rs2$10$ ,\picorv32_core/pcpi_rs2$9$ ,\picorv32_core/pcpi_rs2$8$ ,mem_la_wdata[7:0]}),
    .o(\picorv32_core/alu_lts ));  // ../src/picorv32.v(1195)
  lt_u32_u32 \picorv32_core/lt1  (
    .ci(1'b0),
    .i0({\picorv32_core/pcpi_rs1$31$ ,\picorv32_core/pcpi_rs1$30$ ,\picorv32_core/pcpi_rs1$29$ ,\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$25$ ,\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/pcpi_rs1$23$ ,\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs1$21$ ,\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/pcpi_rs1$19$ ,\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$17$ ,\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/pcpi_rs1$15$ ,\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/pcpi_rs1$11$ ,\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$9$ ,\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/pcpi_rs1$7$ ,\picorv32_core/pcpi_rs1$6$ ,\picorv32_core/pcpi_rs1$5$ ,\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/pcpi_rs1$3$ ,\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .i1({\picorv32_core/pcpi_rs2$31$ ,\picorv32_core/pcpi_rs2$30$ ,\picorv32_core/pcpi_rs2$29$ ,\picorv32_core/pcpi_rs2$28$ ,\picorv32_core/pcpi_rs2$27$ ,\picorv32_core/pcpi_rs2$26$ ,\picorv32_core/pcpi_rs2$25$ ,\picorv32_core/pcpi_rs2$24$ ,\picorv32_core/pcpi_rs2$23$ ,\picorv32_core/pcpi_rs2$22$ ,\picorv32_core/pcpi_rs2$21$ ,\picorv32_core/pcpi_rs2$20$ ,\picorv32_core/pcpi_rs2$19$ ,\picorv32_core/pcpi_rs2$18$ ,\picorv32_core/pcpi_rs2$17$ ,\picorv32_core/pcpi_rs2$16$ ,\picorv32_core/pcpi_rs2$15$ ,\picorv32_core/pcpi_rs2$14$ ,\picorv32_core/pcpi_rs2$13$ ,\picorv32_core/pcpi_rs2$12$ ,\picorv32_core/pcpi_rs2$11$ ,\picorv32_core/pcpi_rs2$10$ ,\picorv32_core/pcpi_rs2$9$ ,\picorv32_core/pcpi_rs2$8$ ,mem_la_wdata[7:0]}),
    .o(\picorv32_core/alu_ltu ));  // ../src/picorv32.v(1196)
  lt_u5_u5 \picorv32_core/lt2  (
    .ci(1'b1),
    .i0(5'b00100),
    .i1(\picorv32_core/reg_sh ),
    .o(\picorv32_core/n554 ));  // ../src/picorv32.v(1773)
  reg_sr_as_w1 \picorv32_core/mem_do_prefetch_reg  (
    .clk(clk),
    .d(\picorv32_core/n505 ),
    .en(\picorv32_core/u617_sel_is_2_o ),
    .reset(\picorv32_core/n747 ),
    .set(1'b0),
    .q(\picorv32_core/mem_do_prefetch ));  // ../src/picorv32.v(1906)
  reg_ar_ss_w1 \picorv32_core/mem_do_rdata_reg  (
    .clk(clk),
    .d(1'b0),
    .en(\picorv32_core/n747 ),
    .reset(1'b0),
    .set(\picorv32_core/n731 ),
    .q(\picorv32_core/mem_do_rdata ));  // ../src/picorv32.v(1906)
  reg_ar_ss_w1 \picorv32_core/mem_do_rinst_reg  (
    .clk(clk),
    .d(\picorv32_core/n749 ),
    .en(1'b1),
    .reset(1'b0),
    .set(\picorv32_core/n728 ),
    .q(\picorv32_core/mem_do_rinst ));  // ../src/picorv32.v(1906)
  reg_ar_ss_w1 \picorv32_core/mem_do_wdata_reg  (
    .clk(clk),
    .d(1'b0),
    .en(\picorv32_core/n747 ),
    .reset(1'b0),
    .set(\picorv32_core/n729 ),
    .q(\picorv32_core/mem_do_wdata ));  // ../src/picorv32.v(1906)
  not \picorv32_core/mem_done_inv  (\picorv32_core/mem_done_neg , \picorv32_core/mem_done );
  not \picorv32_core/mem_la_firstword_inv  (\picorv32_core/mem_la_firstword_neg , \picorv32_core/mem_la_firstword );
  not \picorv32_core/mem_la_read_inv  (\picorv32_core/mem_la_read_neg , \picorv32_core/mem_la_read );
  not \picorv32_core/mem_la_secondword_inv  (\picorv32_core/mem_la_secondword_neg , \picorv32_core/mem_la_secondword );
  reg_sr_as_w1 \picorv32_core/mem_la_secondword_reg  (
    .clk(clk),
    .d(\picorv32_core/mem_la_read ),
    .en(\picorv32_core/mux59_sel_is_5_o ),
    .reset(\picorv32_core/n111 ),
    .set(1'b0),
    .q(\picorv32_core/mem_la_secondword ));  // ../src/picorv32.v(605)
  not \picorv32_core/mem_la_use_prefetched_high_word_inv  (\picorv32_core/mem_la_use_prefetched_high_word_neg , \picorv32_core/mem_la_use_prefetched_high_word );
  not \picorv32_core/mem_rdata_latched[0]_inv  (\picorv32_core/mem_rdata_latched$0$_neg , \picorv32_core/mem_rdata_latched [0]);
  not \picorv32_core/mem_rdata_latched[13]_inv  (\picorv32_core/mem_rdata_latched$13$_neg , \picorv32_core/mem_rdata_latched [13]);
  not \picorv32_core/mem_rdata_latched[14]_inv  (\picorv32_core/mem_rdata_latched$14$_neg , \picorv32_core/mem_rdata_latched [14]);
  not \picorv32_core/mem_rdata_latched[15]_inv  (\picorv32_core/mem_rdata_latched$15$_neg , \picorv32_core/mem_rdata_latched [15]);
  not \picorv32_core/mem_rdata_latched[1]_inv  (\picorv32_core/mem_rdata_latched$1$_neg , \picorv32_core/mem_rdata_latched [1]);
  not \picorv32_core/mem_state[1]_inv  (\picorv32_core/mem_state$1$_neg , \picorv32_core/mem_state [1]);
  reg_sr_as_w1 \picorv32_core/mem_valid_reg  (
    .clk(clk),
    .d(\picorv32_core/n148 ),
    .en(1'b1),
    .reset(\picorv32_core/n111 ),
    .set(1'b0),
    .q(\picorv32_core/mem_valid ));  // ../src/picorv32.v(605)
  not \picorv32_core/mem_wordsize[0]_inv  (\picorv32_core/mem_wordsize$0$_neg , \picorv32_core/mem_wordsize [0]);
  not \picorv32_core/mem_wordsize[1]_inv  (\picorv32_core/mem_wordsize$1$_neg , \picorv32_core/mem_wordsize [1]);
  binary_mux_s1_w1 \picorv32_core/mux0_b10  (
    .i0(\picorv32_core/pcpi_rs1$10$ ),
    .i1(\picorv32_core/n30 [8]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[10]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b11  (
    .i0(\picorv32_core/pcpi_rs1$11$ ),
    .i1(\picorv32_core/n30 [9]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[11]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b12  (
    .i0(\picorv32_core/pcpi_rs1$12$ ),
    .i1(\picorv32_core/n30 [10]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[12]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b13  (
    .i0(\picorv32_core/pcpi_rs1$13$ ),
    .i1(\picorv32_core/n30 [11]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[13]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b14  (
    .i0(\picorv32_core/pcpi_rs1$14$ ),
    .i1(\picorv32_core/n30 [12]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[14]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b15  (
    .i0(\picorv32_core/pcpi_rs1$15$ ),
    .i1(\picorv32_core/n30 [13]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[15]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b16  (
    .i0(\picorv32_core/pcpi_rs1$16$ ),
    .i1(\picorv32_core/n30 [14]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[16]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b17  (
    .i0(\picorv32_core/pcpi_rs1$17$ ),
    .i1(\picorv32_core/n30 [15]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[17]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b18  (
    .i0(\picorv32_core/pcpi_rs1$18$ ),
    .i1(\picorv32_core/n30 [16]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[18]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b19  (
    .i0(\picorv32_core/pcpi_rs1$19$ ),
    .i1(\picorv32_core/n30 [17]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[19]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b2  (
    .i0(\picorv32_core/pcpi_rs1$2$ ),
    .i1(\picorv32_core/n30 [0]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[2]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b20  (
    .i0(\picorv32_core/pcpi_rs1$20$ ),
    .i1(\picorv32_core/n30 [18]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[20]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b21  (
    .i0(\picorv32_core/pcpi_rs1$21$ ),
    .i1(\picorv32_core/n30 [19]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[21]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b22  (
    .i0(\picorv32_core/pcpi_rs1$22$ ),
    .i1(\picorv32_core/n30 [20]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[22]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b23  (
    .i0(\picorv32_core/pcpi_rs1$23$ ),
    .i1(\picorv32_core/n30 [21]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[23]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b24  (
    .i0(\picorv32_core/pcpi_rs1$24$ ),
    .i1(\picorv32_core/n30 [22]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[24]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b25  (
    .i0(\picorv32_core/pcpi_rs1$25$ ),
    .i1(\picorv32_core/n30 [23]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[25]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b26  (
    .i0(\picorv32_core/pcpi_rs1$26$ ),
    .i1(\picorv32_core/n30 [24]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[26]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b27  (
    .i0(\picorv32_core/pcpi_rs1$27$ ),
    .i1(\picorv32_core/n30 [25]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[27]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b28  (
    .i0(\picorv32_core/pcpi_rs1$28$ ),
    .i1(\picorv32_core/n30 [26]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[28]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b29  (
    .i0(\picorv32_core/pcpi_rs1$29$ ),
    .i1(\picorv32_core/n30 [27]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[29]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b3  (
    .i0(\picorv32_core/pcpi_rs1$3$ ),
    .i1(\picorv32_core/n30 [1]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[3]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b30  (
    .i0(\picorv32_core/pcpi_rs1$30$ ),
    .i1(\picorv32_core/n30 [28]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[30]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b31  (
    .i0(\picorv32_core/pcpi_rs1$31$ ),
    .i1(\picorv32_core/n30 [29]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[31]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b4  (
    .i0(\picorv32_core/pcpi_rs1$4$ ),
    .i1(\picorv32_core/n30 [2]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[4]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b5  (
    .i0(\picorv32_core/pcpi_rs1$5$ ),
    .i1(\picorv32_core/n30 [3]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[5]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b6  (
    .i0(\picorv32_core/pcpi_rs1$6$ ),
    .i1(\picorv32_core/n30 [4]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[6]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b7  (
    .i0(\picorv32_core/pcpi_rs1$7$ ),
    .i1(\picorv32_core/n30 [5]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[7]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b8  (
    .i0(\picorv32_core/pcpi_rs1$8$ ),
    .i1(\picorv32_core/n30 [6]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[8]));  // ../src/picorv32.v(346)
  binary_mux_s1_w1 \picorv32_core/mux0_b9  (
    .i0(\picorv32_core/pcpi_rs1$9$ ),
    .i1(\picorv32_core/n30 [7]),
    .sel(\picorv32_core/n0 ),
    .o(mem_la_addr[9]));  // ../src/picorv32.v(346)
  and \picorv32_core/mux100_sel_is_6  (\picorv32_core/mux100_sel_is_6_o , \picorv32_core/mem_rdata_latched$0$_neg , \picorv32_core/mem_rdata_latched [1], \picorv32_core/u247_sel_is_1_o );
  binary_mux_s2_w1 \picorv32_core/mux101  (
    .i0(\picorv32_core/n179 ),
    .i1(\picorv32_core/n213 ),
    .i2(\picorv32_core/n233 ),
    .i3(\picorv32_core/n179 ),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n240 ));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux102  (
    .i0(\picorv32_core/n191 ),
    .i1(\picorv32_core/n177 ),
    .i2(\picorv32_core/n191 ),
    .i3(\picorv32_core/n177 ),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n241 ));  // ../src/picorv32.v(989)
  and \picorv32_core/mux103_sel_is_5  (\picorv32_core/mux103_sel_is_5_o , \picorv32_core/mem_rdata_latched [0], \picorv32_core/mem_rdata_latched$1$_neg , \picorv32_core/mux12_b0_sel_is_3_o );
  and \picorv32_core/mux104_sel_is_5  (\picorv32_core/mux104_sel_is_5_o , \picorv32_core/mem_rdata_latched [0], \picorv32_core/mem_rdata_latched$1$_neg , \picorv32_core/mux81_sel_is_1_o );
  and \picorv32_core/mux105_sel_is_5  (\picorv32_core/mux105_sel_is_5_o , \picorv32_core/mem_rdata_latched [0], \picorv32_core/mem_rdata_latched$1$_neg , \picorv32_core/mux24_b3_sel_is_3_o );
  binary_mux_s1_w1 \picorv32_core/mux106_b0  (
    .i0(\picorv32_core/mem_rdata_latched [7]),
    .i1(\picorv32_core/n235 [0]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n245 [0]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux106_b1  (
    .i0(\picorv32_core/mem_rdata_latched [8]),
    .i1(\picorv32_core/n235 [1]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n245 [1]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux106_b2  (
    .i0(\picorv32_core/mem_rdata_latched [9]),
    .i1(\picorv32_core/n235 [2]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n245 [2]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux106_b3  (
    .i0(\picorv32_core/mem_rdata_latched [10]),
    .i1(\picorv32_core/n235 [3]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n245 [3]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux106_b4  (
    .i0(\picorv32_core/mem_rdata_latched [11]),
    .i1(\picorv32_core/n235 [4]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n245 [4]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux107_b0  (
    .i0(\picorv32_core/mem_rdata_latched [15]),
    .i1(\picorv32_core/n236 [0]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n246 [0]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux107_b1  (
    .i0(\picorv32_core/mem_rdata_latched [16]),
    .i1(\picorv32_core/n236 [1]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n246 [1]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux107_b2  (
    .i0(\picorv32_core/mem_rdata_latched [17]),
    .i1(\picorv32_core/n236 [2]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n246 [2]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux107_b3  (
    .i0(\picorv32_core/mem_rdata_latched [18]),
    .i1(\picorv32_core/n236 [3]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n246 [3]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux107_b4  (
    .i0(\picorv32_core/mem_rdata_latched [19]),
    .i1(\picorv32_core/n236 [4]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n246 [4]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux108_b0  (
    .i0(\picorv32_core/mem_rdata_latched [20]),
    .i1(\picorv32_core/n237 [0]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n247 [0]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux108_b1  (
    .i0(\picorv32_core/mem_rdata_latched [21]),
    .i1(\picorv32_core/n237 [1]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n247 [1]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux108_b2  (
    .i0(\picorv32_core/mem_rdata_latched [22]),
    .i1(\picorv32_core/n237 [2]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n247 [2]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux108_b3  (
    .i0(\picorv32_core/mem_rdata_latched [23]),
    .i1(\picorv32_core/n237 [3]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n247 [3]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux108_b4  (
    .i0(\picorv32_core/mem_rdata_latched [24]),
    .i1(\picorv32_core/n237 [4]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n247 [4]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux10_b10  (
    .i0(\picorv32_core/mem_rdata_q [10]),
    .i1(\picorv32_core/mem_rdata_latched [10]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [10]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b11  (
    .i0(\picorv32_core/mem_rdata_q [11]),
    .i1(\picorv32_core/mem_rdata_latched [11]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [11]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b12  (
    .i0(\picorv32_core/mem_rdata_q [12]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [12]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b13  (
    .i0(\picorv32_core/mem_rdata_q [13]),
    .i1(\picorv32_core/mem_rdata_latched [13]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [13]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b14  (
    .i0(\picorv32_core/mem_rdata_q [14]),
    .i1(\picorv32_core/mem_rdata_latched [14]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [14]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b15  (
    .i0(\picorv32_core/mem_rdata_q [15]),
    .i1(\picorv32_core/mem_rdata_latched [15]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [15]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b16  (
    .i0(\picorv32_core/mem_rdata_q [16]),
    .i1(\picorv32_core/mem_rdata_latched [16]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [16]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b17  (
    .i0(\picorv32_core/mem_rdata_q [17]),
    .i1(\picorv32_core/mem_rdata_latched [17]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [17]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b18  (
    .i0(\picorv32_core/mem_rdata_q [18]),
    .i1(\picorv32_core/mem_rdata_latched [18]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [18]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b19  (
    .i0(\picorv32_core/mem_rdata_q [19]),
    .i1(\picorv32_core/mem_rdata_latched [19]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [19]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b20  (
    .i0(\picorv32_core/mem_rdata_q [20]),
    .i1(\picorv32_core/mem_rdata_latched [20]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [20]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b21  (
    .i0(\picorv32_core/mem_rdata_q [21]),
    .i1(\picorv32_core/mem_rdata_latched [21]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [21]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b22  (
    .i0(\picorv32_core/mem_rdata_q [22]),
    .i1(\picorv32_core/mem_rdata_latched [22]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [22]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b23  (
    .i0(\picorv32_core/mem_rdata_q [23]),
    .i1(\picorv32_core/mem_rdata_latched [23]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [23]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b24  (
    .i0(\picorv32_core/mem_rdata_q [24]),
    .i1(\picorv32_core/mem_rdata_latched [24]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [24]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b25  (
    .i0(\picorv32_core/mem_rdata_q [25]),
    .i1(\picorv32_core/mem_rdata_latched [25]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [25]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b26  (
    .i0(\picorv32_core/mem_rdata_q [26]),
    .i1(\picorv32_core/mem_rdata_latched [26]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [26]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b27  (
    .i0(\picorv32_core/mem_rdata_q [27]),
    .i1(\picorv32_core/mem_rdata_latched [27]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [27]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b28  (
    .i0(\picorv32_core/mem_rdata_q [28]),
    .i1(\picorv32_core/mem_rdata_latched [28]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [28]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b29  (
    .i0(\picorv32_core/mem_rdata_q [29]),
    .i1(\picorv32_core/mem_rdata_latched [29]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [29]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b30  (
    .i0(\picorv32_core/mem_rdata_q [30]),
    .i1(\picorv32_core/mem_rdata_latched [30]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [30]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b31  (
    .i0(\picorv32_core/mem_rdata_q [31]),
    .i1(\picorv32_core/mem_rdata_latched [31]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [31]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b7  (
    .i0(\picorv32_core/mem_rdata_q [7]),
    .i1(\picorv32_core/mem_rdata_latched [7]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [7]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b8  (
    .i0(\picorv32_core/mem_rdata_q [8]),
    .i1(\picorv32_core/mem_rdata_latched [8]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [8]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux10_b9  (
    .i0(\picorv32_core/mem_rdata_q [9]),
    .i1(\picorv32_core/mem_rdata_latched [9]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n42 [9]));  // ../src/picorv32.v(398)
  binary_mux_s1_w1 \picorv32_core/mux115_b1  (
    .i0(\picorv32_core/reg_next_pc [1]),
    .i1(\picorv32_core/reg_out [1]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [1]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b10  (
    .i0(\picorv32_core/reg_next_pc [10]),
    .i1(\picorv32_core/reg_out [10]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [10]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b11  (
    .i0(\picorv32_core/reg_next_pc [11]),
    .i1(\picorv32_core/reg_out [11]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [11]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b12  (
    .i0(\picorv32_core/reg_next_pc [12]),
    .i1(\picorv32_core/reg_out [12]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [12]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b13  (
    .i0(\picorv32_core/reg_next_pc [13]),
    .i1(\picorv32_core/reg_out [13]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [13]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b14  (
    .i0(\picorv32_core/reg_next_pc [14]),
    .i1(\picorv32_core/reg_out [14]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [14]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b15  (
    .i0(\picorv32_core/reg_next_pc [15]),
    .i1(\picorv32_core/reg_out [15]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [15]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b16  (
    .i0(\picorv32_core/reg_next_pc [16]),
    .i1(\picorv32_core/reg_out [16]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [16]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b17  (
    .i0(\picorv32_core/reg_next_pc [17]),
    .i1(\picorv32_core/reg_out [17]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [17]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b18  (
    .i0(\picorv32_core/reg_next_pc [18]),
    .i1(\picorv32_core/reg_out [18]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [18]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b19  (
    .i0(\picorv32_core/reg_next_pc [19]),
    .i1(\picorv32_core/reg_out [19]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [19]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b2  (
    .i0(\picorv32_core/reg_next_pc [2]),
    .i1(\picorv32_core/reg_out [2]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [2]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b20  (
    .i0(\picorv32_core/reg_next_pc [20]),
    .i1(\picorv32_core/reg_out [20]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [20]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b21  (
    .i0(\picorv32_core/reg_next_pc [21]),
    .i1(\picorv32_core/reg_out [21]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [21]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b22  (
    .i0(\picorv32_core/reg_next_pc [22]),
    .i1(\picorv32_core/reg_out [22]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [22]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b23  (
    .i0(\picorv32_core/reg_next_pc [23]),
    .i1(\picorv32_core/reg_out [23]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [23]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b24  (
    .i0(\picorv32_core/reg_next_pc [24]),
    .i1(\picorv32_core/reg_out [24]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [24]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b25  (
    .i0(\picorv32_core/reg_next_pc [25]),
    .i1(\picorv32_core/reg_out [25]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [25]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b26  (
    .i0(\picorv32_core/reg_next_pc [26]),
    .i1(\picorv32_core/reg_out [26]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [26]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b27  (
    .i0(\picorv32_core/reg_next_pc [27]),
    .i1(\picorv32_core/reg_out [27]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [27]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b28  (
    .i0(\picorv32_core/reg_next_pc [28]),
    .i1(\picorv32_core/reg_out [28]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [28]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b29  (
    .i0(\picorv32_core/reg_next_pc [29]),
    .i1(\picorv32_core/reg_out [29]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [29]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b3  (
    .i0(\picorv32_core/reg_next_pc [3]),
    .i1(\picorv32_core/reg_out [3]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [3]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b30  (
    .i0(\picorv32_core/reg_next_pc [30]),
    .i1(\picorv32_core/reg_out [30]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [30]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b31  (
    .i0(\picorv32_core/reg_next_pc [31]),
    .i1(\picorv32_core/reg_out [31]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [31]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b4  (
    .i0(\picorv32_core/reg_next_pc [4]),
    .i1(\picorv32_core/reg_out [4]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [4]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b5  (
    .i0(\picorv32_core/reg_next_pc [5]),
    .i1(\picorv32_core/reg_out [5]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [5]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b6  (
    .i0(\picorv32_core/reg_next_pc [6]),
    .i1(\picorv32_core/reg_out [6]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [6]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b7  (
    .i0(\picorv32_core/reg_next_pc [7]),
    .i1(\picorv32_core/reg_out [7]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [7]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b8  (
    .i0(\picorv32_core/reg_next_pc [8]),
    .i1(\picorv32_core/reg_out [8]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [8]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux115_b9  (
    .i0(\picorv32_core/reg_next_pc [9]),
    .i1(\picorv32_core/reg_out [9]),
    .sel(\picorv32_core/n432 ),
    .o(\picorv32_core/next_pc [9]));  // ../src/picorv32.v(1166)
  binary_mux_s1_w1 \picorv32_core/mux116_b0  (
    .i0(\picorv32_core/n434 [0]),
    .i1(\picorv32_core/n433 [0]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [0]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b1  (
    .i0(\picorv32_core/n434 [1]),
    .i1(\picorv32_core/n433 [1]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [1]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b10  (
    .i0(\picorv32_core/n434 [10]),
    .i1(\picorv32_core/n433 [10]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [10]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b11  (
    .i0(\picorv32_core/n434 [11]),
    .i1(\picorv32_core/n433 [11]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [11]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b12  (
    .i0(\picorv32_core/n434 [12]),
    .i1(\picorv32_core/n433 [12]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [12]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b13  (
    .i0(\picorv32_core/n434 [13]),
    .i1(\picorv32_core/n433 [13]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [13]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b14  (
    .i0(\picorv32_core/n434 [14]),
    .i1(\picorv32_core/n433 [14]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [14]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b15  (
    .i0(\picorv32_core/n434 [15]),
    .i1(\picorv32_core/n433 [15]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [15]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b16  (
    .i0(\picorv32_core/n434 [16]),
    .i1(\picorv32_core/n433 [16]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [16]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b17  (
    .i0(\picorv32_core/n434 [17]),
    .i1(\picorv32_core/n433 [17]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [17]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b18  (
    .i0(\picorv32_core/n434 [18]),
    .i1(\picorv32_core/n433 [18]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [18]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b19  (
    .i0(\picorv32_core/n434 [19]),
    .i1(\picorv32_core/n433 [19]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [19]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b2  (
    .i0(\picorv32_core/n434 [2]),
    .i1(\picorv32_core/n433 [2]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [2]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b20  (
    .i0(\picorv32_core/n434 [20]),
    .i1(\picorv32_core/n433 [20]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [20]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b21  (
    .i0(\picorv32_core/n434 [21]),
    .i1(\picorv32_core/n433 [21]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [21]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b22  (
    .i0(\picorv32_core/n434 [22]),
    .i1(\picorv32_core/n433 [22]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [22]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b23  (
    .i0(\picorv32_core/n434 [23]),
    .i1(\picorv32_core/n433 [23]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [23]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b24  (
    .i0(\picorv32_core/n434 [24]),
    .i1(\picorv32_core/n433 [24]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [24]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b25  (
    .i0(\picorv32_core/n434 [25]),
    .i1(\picorv32_core/n433 [25]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [25]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b26  (
    .i0(\picorv32_core/n434 [26]),
    .i1(\picorv32_core/n433 [26]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [26]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b27  (
    .i0(\picorv32_core/n434 [27]),
    .i1(\picorv32_core/n433 [27]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [27]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b28  (
    .i0(\picorv32_core/n434 [28]),
    .i1(\picorv32_core/n433 [28]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [28]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b29  (
    .i0(\picorv32_core/n434 [29]),
    .i1(\picorv32_core/n433 [29]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [29]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b3  (
    .i0(\picorv32_core/n434 [3]),
    .i1(\picorv32_core/n433 [3]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [3]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b30  (
    .i0(\picorv32_core/n434 [30]),
    .i1(\picorv32_core/n433 [30]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [30]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b31  (
    .i0(\picorv32_core/n434 [31]),
    .i1(\picorv32_core/n433 [31]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [31]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b4  (
    .i0(\picorv32_core/n434 [4]),
    .i1(\picorv32_core/n433 [4]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [4]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b5  (
    .i0(\picorv32_core/n434 [5]),
    .i1(\picorv32_core/n433 [5]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [5]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b6  (
    .i0(\picorv32_core/n434 [6]),
    .i1(\picorv32_core/n433 [6]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [6]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b7  (
    .i0(\picorv32_core/n434 [7]),
    .i1(\picorv32_core/n433 [7]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [7]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b8  (
    .i0(\picorv32_core/n434 [8]),
    .i1(\picorv32_core/n433 [8]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [8]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux116_b9  (
    .i0(\picorv32_core/n434 [9]),
    .i1(\picorv32_core/n433 [9]),
    .sel(\picorv32_core/instr_sub ),
    .o(\picorv32_core/alu_add_sub [9]));  // ../src/picorv32.v(1193)
  binary_mux_s1_w1 \picorv32_core/mux117_b0  (
    .i0(\picorv32_core/reg_out [0]),
    .i1(\picorv32_core/alu_out_q [0]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [0]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b1  (
    .i0(\picorv32_core/reg_out [1]),
    .i1(\picorv32_core/alu_out_q [1]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [1]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b10  (
    .i0(\picorv32_core/reg_out [10]),
    .i1(\picorv32_core/alu_out_q [10]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [10]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b11  (
    .i0(\picorv32_core/reg_out [11]),
    .i1(\picorv32_core/alu_out_q [11]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [11]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b12  (
    .i0(\picorv32_core/reg_out [12]),
    .i1(\picorv32_core/alu_out_q [12]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [12]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b13  (
    .i0(\picorv32_core/reg_out [13]),
    .i1(\picorv32_core/alu_out_q [13]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [13]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b14  (
    .i0(\picorv32_core/reg_out [14]),
    .i1(\picorv32_core/alu_out_q [14]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [14]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b15  (
    .i0(\picorv32_core/reg_out [15]),
    .i1(\picorv32_core/alu_out_q [15]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [15]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b16  (
    .i0(\picorv32_core/reg_out [16]),
    .i1(\picorv32_core/alu_out_q [16]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [16]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b17  (
    .i0(\picorv32_core/reg_out [17]),
    .i1(\picorv32_core/alu_out_q [17]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [17]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b18  (
    .i0(\picorv32_core/reg_out [18]),
    .i1(\picorv32_core/alu_out_q [18]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [18]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b19  (
    .i0(\picorv32_core/reg_out [19]),
    .i1(\picorv32_core/alu_out_q [19]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [19]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b2  (
    .i0(\picorv32_core/reg_out [2]),
    .i1(\picorv32_core/alu_out_q [2]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [2]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b20  (
    .i0(\picorv32_core/reg_out [20]),
    .i1(\picorv32_core/alu_out_q [20]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [20]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b21  (
    .i0(\picorv32_core/reg_out [21]),
    .i1(\picorv32_core/alu_out_q [21]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [21]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b22  (
    .i0(\picorv32_core/reg_out [22]),
    .i1(\picorv32_core/alu_out_q [22]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [22]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b23  (
    .i0(\picorv32_core/reg_out [23]),
    .i1(\picorv32_core/alu_out_q [23]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [23]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b24  (
    .i0(\picorv32_core/reg_out [24]),
    .i1(\picorv32_core/alu_out_q [24]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [24]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b25  (
    .i0(\picorv32_core/reg_out [25]),
    .i1(\picorv32_core/alu_out_q [25]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [25]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b26  (
    .i0(\picorv32_core/reg_out [26]),
    .i1(\picorv32_core/alu_out_q [26]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [26]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b27  (
    .i0(\picorv32_core/reg_out [27]),
    .i1(\picorv32_core/alu_out_q [27]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [27]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b28  (
    .i0(\picorv32_core/reg_out [28]),
    .i1(\picorv32_core/alu_out_q [28]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [28]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b29  (
    .i0(\picorv32_core/reg_out [29]),
    .i1(\picorv32_core/alu_out_q [29]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [29]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b3  (
    .i0(\picorv32_core/reg_out [3]),
    .i1(\picorv32_core/alu_out_q [3]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [3]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b30  (
    .i0(\picorv32_core/reg_out [30]),
    .i1(\picorv32_core/alu_out_q [30]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [30]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b31  (
    .i0(\picorv32_core/reg_out [31]),
    .i1(\picorv32_core/alu_out_q [31]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [31]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b4  (
    .i0(\picorv32_core/reg_out [4]),
    .i1(\picorv32_core/alu_out_q [4]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [4]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b5  (
    .i0(\picorv32_core/reg_out [5]),
    .i1(\picorv32_core/alu_out_q [5]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [5]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b6  (
    .i0(\picorv32_core/reg_out [6]),
    .i1(\picorv32_core/alu_out_q [6]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [6]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b7  (
    .i0(\picorv32_core/reg_out [7]),
    .i1(\picorv32_core/alu_out_q [7]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [7]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b8  (
    .i0(\picorv32_core/reg_out [8]),
    .i1(\picorv32_core/alu_out_q [8]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [8]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux117_b9  (
    .i0(\picorv32_core/reg_out [9]),
    .i1(\picorv32_core/alu_out_q [9]),
    .sel(\picorv32_core/latched_stalu ),
    .o(\picorv32_core/n453 [9]));  // ../src/picorv32.v(1274)
  binary_mux_s1_w1 \picorv32_core/mux118_b0  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [0]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [0]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b1  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [1]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [1]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b10  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [10]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [10]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b11  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [11]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [11]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b12  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [12]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [12]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b13  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [13]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [13]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b14  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [14]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [14]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b15  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [15]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [15]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b16  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [16]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [16]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b17  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [17]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [17]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b18  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [18]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [18]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b19  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [19]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [19]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b2  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [2]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [2]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b20  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [20]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [20]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b21  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [21]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [21]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b22  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [22]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [22]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b23  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [23]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [23]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b24  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [24]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [24]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b25  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [25]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [25]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b26  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [26]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [26]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b27  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [27]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [27]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b28  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [28]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [28]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b29  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [29]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [29]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b3  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [3]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [3]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b30  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [30]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [30]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b31  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [31]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [31]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b4  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [4]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [4]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b5  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [5]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [5]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b6  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [6]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [6]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b7  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [7]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [7]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b8  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [8]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [8]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux118_b9  (
    .i0(1'bx),
    .i1(\picorv32_core/n455 [9]),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_wrdata [9]));  // ../src/picorv32.v(1286)
  binary_mux_s1_w1 \picorv32_core/mux119_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [0]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [0]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [1]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [1]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b10  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [10]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [10]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b11  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [11]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [11]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b12  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [12]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [12]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b13  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [13]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [13]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b14  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [14]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [14]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b15  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [15]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [15]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b16  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [16]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [16]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b17  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [17]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [17]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b18  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [18]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [18]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b19  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [19]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [19]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b2  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [2]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [2]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b20  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [20]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [20]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b21  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [21]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [21]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b22  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [22]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [22]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b23  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [23]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [23]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b24  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [24]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [24]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b25  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [25]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [25]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b26  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [26]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [26]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b27  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [27]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [27]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b28  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [28]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [28]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b29  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [29]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [29]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b3  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [3]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [3]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b30  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [30]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [30]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b31  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [31]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [31]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b4  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [4]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [4]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b5  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [5]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [5]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b6  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [6]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [6]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b7  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [7]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [7]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b8  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [8]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [8]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux119_b9  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs1_z [9]),
    .sel(\picorv32_core/n457 ),
    .o(\picorv32_core/cpuregs_rs1 [9]));  // ../src/picorv32.v(1328)
  binary_mux_s1_w1 \picorv32_core/mux11_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [2]),
    .sel(\picorv32_core/n188 ),
    .o(\picorv32_core/n189 [0]));  // ../src/picorv32.v(882)
  binary_mux_s1_w1 \picorv32_core/mux11_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [3]),
    .sel(\picorv32_core/n188 ),
    .o(\picorv32_core/n189 [1]));  // ../src/picorv32.v(882)
  binary_mux_s1_w1 \picorv32_core/mux11_b2  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [4]),
    .sel(\picorv32_core/n188 ),
    .o(\picorv32_core/n189 [2]));  // ../src/picorv32.v(882)
  binary_mux_s1_w1 \picorv32_core/mux120_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [0]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [0]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [1]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [1]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b10  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [10]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [10]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b11  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [11]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [11]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b12  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [12]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [12]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b13  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [13]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [13]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b14  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [14]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [14]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b15  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [15]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [15]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b16  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [16]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [16]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b17  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [17]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [17]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b18  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [18]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [18]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b19  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [19]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [19]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b2  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [2]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [2]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b20  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [20]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [20]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b21  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [21]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [21]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b22  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [22]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [22]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b23  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [23]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [23]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b24  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [24]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [24]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b25  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [25]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [25]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b26  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [26]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [26]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b27  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [27]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [27]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b28  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [28]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [28]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b29  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [29]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [29]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b3  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [3]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [3]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b30  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [30]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [30]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b31  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [31]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [31]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b4  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [4]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [4]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b5  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [5]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [5]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b6  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [6]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [6]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b7  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [7]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [7]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b8  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [8]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [8]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux120_b9  (
    .i0(1'b0),
    .i1(\picorv32_core/cpuregs_rs2_z [9]),
    .sel(\picorv32_core/n458 ),
    .o(\picorv32_core/cpuregs_rs2 [9]));  // ../src/picorv32.v(1329)
  binary_mux_s1_w1 \picorv32_core/mux123_b0  (
    .i0(\picorv32_core/n502 [0]),
    .i1(\picorv32_core/n504 [0]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [0]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b1  (
    .i0(\picorv32_core/n502 [1]),
    .i1(\picorv32_core/n504 [1]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [1]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b10  (
    .i0(\picorv32_core/n502 [10]),
    .i1(\picorv32_core/n504 [10]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [10]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b11  (
    .i0(\picorv32_core/n502 [11]),
    .i1(\picorv32_core/n504 [11]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [11]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b12  (
    .i0(\picorv32_core/n502 [12]),
    .i1(\picorv32_core/n504 [12]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [12]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b13  (
    .i0(\picorv32_core/n502 [13]),
    .i1(\picorv32_core/n504 [13]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [13]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b14  (
    .i0(\picorv32_core/n502 [14]),
    .i1(\picorv32_core/n504 [14]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [14]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b15  (
    .i0(\picorv32_core/n502 [15]),
    .i1(\picorv32_core/n504 [15]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [15]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b16  (
    .i0(\picorv32_core/n502 [16]),
    .i1(\picorv32_core/n504 [16]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [16]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b17  (
    .i0(\picorv32_core/n502 [17]),
    .i1(\picorv32_core/n504 [17]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [17]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b18  (
    .i0(\picorv32_core/n502 [18]),
    .i1(\picorv32_core/n504 [18]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [18]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b19  (
    .i0(\picorv32_core/n502 [19]),
    .i1(\picorv32_core/n504 [19]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [19]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b2  (
    .i0(\picorv32_core/n502 [2]),
    .i1(\picorv32_core/n504 [2]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [2]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b20  (
    .i0(\picorv32_core/n502 [20]),
    .i1(\picorv32_core/n504 [20]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [20]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b21  (
    .i0(\picorv32_core/n502 [21]),
    .i1(\picorv32_core/n504 [21]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [21]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b22  (
    .i0(\picorv32_core/n502 [22]),
    .i1(\picorv32_core/n504 [22]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [22]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b23  (
    .i0(\picorv32_core/n502 [23]),
    .i1(\picorv32_core/n504 [23]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [23]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b24  (
    .i0(\picorv32_core/n502 [24]),
    .i1(\picorv32_core/n504 [24]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [24]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b25  (
    .i0(\picorv32_core/n502 [25]),
    .i1(\picorv32_core/n504 [25]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [25]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b26  (
    .i0(\picorv32_core/n502 [26]),
    .i1(\picorv32_core/n504 [26]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [26]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b27  (
    .i0(\picorv32_core/n502 [27]),
    .i1(\picorv32_core/n504 [27]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [27]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b28  (
    .i0(\picorv32_core/n502 [28]),
    .i1(\picorv32_core/n504 [28]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [28]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b29  (
    .i0(\picorv32_core/n502 [29]),
    .i1(\picorv32_core/n504 [29]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [29]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b3  (
    .i0(\picorv32_core/n502 [3]),
    .i1(\picorv32_core/n504 [3]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [3]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b30  (
    .i0(\picorv32_core/n502 [30]),
    .i1(\picorv32_core/n504 [30]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [30]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b31  (
    .i0(\picorv32_core/n502 [31]),
    .i1(\picorv32_core/n504 [31]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [31]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b4  (
    .i0(\picorv32_core/n502 [4]),
    .i1(\picorv32_core/n504 [4]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [4]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b5  (
    .i0(\picorv32_core/n502 [5]),
    .i1(\picorv32_core/n504 [5]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [5]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b6  (
    .i0(\picorv32_core/n502 [6]),
    .i1(\picorv32_core/n504 [6]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [6]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b7  (
    .i0(\picorv32_core/n502 [7]),
    .i1(\picorv32_core/n504 [7]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [7]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b8  (
    .i0(\picorv32_core/n502 [8]),
    .i1(\picorv32_core/n504 [8]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [8]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux123_b9  (
    .i0(\picorv32_core/n502 [9]),
    .i1(\picorv32_core/n504 [9]),
    .sel(\picorv32_core/instr_jal ),
    .o(\picorv32_core/n508 [9]));  // ../src/picorv32.v(1513)
  binary_mux_s1_w1 \picorv32_core/mux125_b0  (
    .i0(\picorv32_core/n500 [0]),
    .i1(\picorv32_core/n508 [0]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [0]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b1  (
    .i0(\picorv32_core/n500 [1]),
    .i1(\picorv32_core/n508 [1]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [1]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b10  (
    .i0(\picorv32_core/n500 [10]),
    .i1(\picorv32_core/n508 [10]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [10]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b11  (
    .i0(\picorv32_core/n500 [11]),
    .i1(\picorv32_core/n508 [11]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [11]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b12  (
    .i0(\picorv32_core/n500 [12]),
    .i1(\picorv32_core/n508 [12]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [12]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b13  (
    .i0(\picorv32_core/n500 [13]),
    .i1(\picorv32_core/n508 [13]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [13]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b14  (
    .i0(\picorv32_core/n500 [14]),
    .i1(\picorv32_core/n508 [14]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [14]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b15  (
    .i0(\picorv32_core/n500 [15]),
    .i1(\picorv32_core/n508 [15]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [15]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b16  (
    .i0(\picorv32_core/n500 [16]),
    .i1(\picorv32_core/n508 [16]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [16]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b17  (
    .i0(\picorv32_core/n500 [17]),
    .i1(\picorv32_core/n508 [17]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [17]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b18  (
    .i0(\picorv32_core/n500 [18]),
    .i1(\picorv32_core/n508 [18]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [18]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b19  (
    .i0(\picorv32_core/n500 [19]),
    .i1(\picorv32_core/n508 [19]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [19]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b2  (
    .i0(\picorv32_core/n500 [2]),
    .i1(\picorv32_core/n508 [2]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [2]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b20  (
    .i0(\picorv32_core/n500 [20]),
    .i1(\picorv32_core/n508 [20]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [20]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b21  (
    .i0(\picorv32_core/n500 [21]),
    .i1(\picorv32_core/n508 [21]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [21]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b22  (
    .i0(\picorv32_core/n500 [22]),
    .i1(\picorv32_core/n508 [22]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [22]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b23  (
    .i0(\picorv32_core/n500 [23]),
    .i1(\picorv32_core/n508 [23]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [23]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b24  (
    .i0(\picorv32_core/n500 [24]),
    .i1(\picorv32_core/n508 [24]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [24]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b25  (
    .i0(\picorv32_core/n500 [25]),
    .i1(\picorv32_core/n508 [25]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [25]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b26  (
    .i0(\picorv32_core/n500 [26]),
    .i1(\picorv32_core/n508 [26]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [26]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b27  (
    .i0(\picorv32_core/n500 [27]),
    .i1(\picorv32_core/n508 [27]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [27]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b28  (
    .i0(\picorv32_core/n500 [28]),
    .i1(\picorv32_core/n508 [28]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [28]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b29  (
    .i0(\picorv32_core/n500 [29]),
    .i1(\picorv32_core/n508 [29]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [29]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b3  (
    .i0(\picorv32_core/n500 [3]),
    .i1(\picorv32_core/n508 [3]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [3]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b30  (
    .i0(\picorv32_core/n500 [30]),
    .i1(\picorv32_core/n508 [30]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [30]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b31  (
    .i0(\picorv32_core/n500 [31]),
    .i1(\picorv32_core/n508 [31]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [31]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b4  (
    .i0(\picorv32_core/n500 [4]),
    .i1(\picorv32_core/n508 [4]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [4]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b5  (
    .i0(\picorv32_core/n500 [5]),
    .i1(\picorv32_core/n508 [5]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [5]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b6  (
    .i0(\picorv32_core/n500 [6]),
    .i1(\picorv32_core/n508 [6]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [6]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b7  (
    .i0(\picorv32_core/n500 [7]),
    .i1(\picorv32_core/n508 [7]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [7]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b8  (
    .i0(\picorv32_core/n500 [8]),
    .i1(\picorv32_core/n508 [8]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [8]));  // ../src/picorv32.v(1514)
  binary_mux_s1_w1 \picorv32_core/mux125_b9  (
    .i0(\picorv32_core/n500 [9]),
    .i1(\picorv32_core/n508 [9]),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n511 [9]));  // ../src/picorv32.v(1514)
  AL_MUX \picorv32_core/mux127_b0  (
    .i0(\picorv32_core/cpu_state [0]),
    .i1(1'b0),
    .sel(\picorv32_core/mux127_b0_sel_is_1_o ),
    .o(\picorv32_core/n516 [0]));
  and \picorv32_core/mux127_b0_sel_is_1  (\picorv32_core/mux127_b0_sel_is_1_o , \picorv32_core/decoder_trigger , \picorv32_core/instr_jal_neg );
  AL_MUX \picorv32_core/mux127_b1  (
    .i0(\picorv32_core/cpu_state [1]),
    .i1(1'b0),
    .sel(\picorv32_core/mux127_b0_sel_is_1_o ),
    .o(\picorv32_core/n516 [1]));
  AL_MUX \picorv32_core/mux127_b2  (
    .i0(\picorv32_core/cpu_state [2]),
    .i1(1'b0),
    .sel(\picorv32_core/mux127_b0_sel_is_1_o ),
    .o(\picorv32_core/n516 [2]));
  AL_MUX \picorv32_core/mux127_b3  (
    .i0(\picorv32_core/cpu_state [3]),
    .i1(1'b0),
    .sel(\picorv32_core/mux127_b0_sel_is_1_o ),
    .o(\picorv32_core/n516 [3]));
  AL_MUX \picorv32_core/mux127_b4  (
    .i0(\picorv32_core/cpu_state [4]),
    .i1(1'b0),
    .sel(\picorv32_core/mux127_b0_sel_is_1_o ),
    .o(\picorv32_core/n516 [4]));
  AL_MUX \picorv32_core/mux127_b5  (
    .i0(\picorv32_core/cpu_state [5]),
    .i1(1'b1),
    .sel(\picorv32_core/mux127_b0_sel_is_1_o ),
    .o(\picorv32_core/n516 [5]));
  AL_MUX \picorv32_core/mux127_b6  (
    .i0(\picorv32_core/cpu_state [6]),
    .i1(1'b0),
    .sel(\picorv32_core/mux127_b0_sel_is_1_o ),
    .o(\picorv32_core/n516 [6]));
  AL_MUX \picorv32_core/mux127_b7  (
    .i0(\picorv32_core/cpu_state [7]),
    .i1(1'b0),
    .sel(\picorv32_core/mux127_b0_sel_is_1_o ),
    .o(\picorv32_core/n516 [7]));
  binary_mux_s1_w1 \picorv32_core/mux128_b0  (
    .i0(\picorv32_core/reg_pc [0]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [0]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b1  (
    .i0(\picorv32_core/reg_pc [1]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [1]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b10  (
    .i0(\picorv32_core/reg_pc [10]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [10]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b11  (
    .i0(\picorv32_core/reg_pc [11]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [11]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b12  (
    .i0(\picorv32_core/reg_pc [12]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [12]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b13  (
    .i0(\picorv32_core/reg_pc [13]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [13]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b14  (
    .i0(\picorv32_core/reg_pc [14]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [14]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b15  (
    .i0(\picorv32_core/reg_pc [15]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [15]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b16  (
    .i0(\picorv32_core/reg_pc [16]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [16]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b17  (
    .i0(\picorv32_core/reg_pc [17]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [17]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b18  (
    .i0(\picorv32_core/reg_pc [18]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [18]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b19  (
    .i0(\picorv32_core/reg_pc [19]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [19]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b2  (
    .i0(\picorv32_core/reg_pc [2]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [2]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b20  (
    .i0(\picorv32_core/reg_pc [20]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [20]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b21  (
    .i0(\picorv32_core/reg_pc [21]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [21]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b22  (
    .i0(\picorv32_core/reg_pc [22]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [22]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b23  (
    .i0(\picorv32_core/reg_pc [23]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [23]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b24  (
    .i0(\picorv32_core/reg_pc [24]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [24]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b25  (
    .i0(\picorv32_core/reg_pc [25]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [25]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b26  (
    .i0(\picorv32_core/reg_pc [26]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [26]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b27  (
    .i0(\picorv32_core/reg_pc [27]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [27]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b28  (
    .i0(\picorv32_core/reg_pc [28]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [28]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b29  (
    .i0(\picorv32_core/reg_pc [29]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [29]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b3  (
    .i0(\picorv32_core/reg_pc [3]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [3]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b30  (
    .i0(\picorv32_core/reg_pc [30]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [30]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b31  (
    .i0(\picorv32_core/reg_pc [31]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [31]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b4  (
    .i0(\picorv32_core/reg_pc [4]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [4]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b5  (
    .i0(\picorv32_core/reg_pc [5]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [5]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b6  (
    .i0(\picorv32_core/reg_pc [6]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [6]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b7  (
    .i0(\picorv32_core/reg_pc [7]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [7]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b8  (
    .i0(\picorv32_core/reg_pc [8]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [8]));  // ../src/picorv32.v(1580)
  binary_mux_s1_w1 \picorv32_core/mux128_b9  (
    .i0(\picorv32_core/reg_pc [9]),
    .i1(1'b0),
    .sel(\picorv32_core/instr_lui ),
    .o(\picorv32_core/n518 [9]));  // ../src/picorv32.v(1580)
  AL_MUX \picorv32_core/mux12_b0  (
    .i0(\picorv32_core/n42 [7]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/mux12_b0_sel_is_3_o ),
    .o(\picorv32_core/n71 [0]));
  and \picorv32_core/mux12_b0_sel_is_3  (\picorv32_core/mux12_b0_sel_is_3_o , \picorv32_core/mem_rdata_latched [14], \picorv32_core/mem_rdata_latched [15]);
  AL_MUX \picorv32_core/mux12_b1  (
    .i0(\picorv32_core/n42 [8]),
    .i1(\picorv32_core/mem_rdata_latched [3]),
    .sel(\picorv32_core/mux12_b0_sel_is_3_o ),
    .o(\picorv32_core/n71 [1]));
  AL_MUX \picorv32_core/mux12_b2  (
    .i0(\picorv32_core/n42 [9]),
    .i1(\picorv32_core/mem_rdata_latched [4]),
    .sel(\picorv32_core/mux12_b0_sel_is_3_o ),
    .o(\picorv32_core/n71 [2]));
  AL_MUX \picorv32_core/mux12_b3  (
    .i0(\picorv32_core/n42 [10]),
    .i1(\picorv32_core/mem_rdata_latched [10]),
    .sel(\picorv32_core/mux12_b0_sel_is_3_o ),
    .o(\picorv32_core/n71 [3]));
  AL_MUX \picorv32_core/mux12_b4  (
    .i0(\picorv32_core/n42 [11]),
    .i1(\picorv32_core/mem_rdata_latched [11]),
    .sel(\picorv32_core/mux12_b0_sel_is_3_o ),
    .o(\picorv32_core/n71 [4]));
  binary_mux_s1_w1 \picorv32_core/mux130_b0  (
    .i0(\picorv32_core/latched_rd [0]),
    .i1(1'b0),
    .sel(\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ),
    .o(\picorv32_core/n546 [0]));  // ../src/picorv32.v(1764)
  binary_mux_s1_w1 \picorv32_core/mux130_b1  (
    .i0(\picorv32_core/latched_rd [1]),
    .i1(1'b0),
    .sel(\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ),
    .o(\picorv32_core/n546 [1]));  // ../src/picorv32.v(1764)
  binary_mux_s1_w1 \picorv32_core/mux130_b2  (
    .i0(\picorv32_core/latched_rd [2]),
    .i1(1'b0),
    .sel(\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ),
    .o(\picorv32_core/n546 [2]));  // ../src/picorv32.v(1764)
  binary_mux_s1_w1 \picorv32_core/mux130_b3  (
    .i0(\picorv32_core/latched_rd [3]),
    .i1(1'b0),
    .sel(\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ),
    .o(\picorv32_core/n546 [3]));  // ../src/picorv32.v(1764)
  binary_mux_s1_w1 \picorv32_core/mux130_b4  (
    .i0(\picorv32_core/latched_rd [4]),
    .i1(1'b0),
    .sel(\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ),
    .o(\picorv32_core/n546 [4]));  // ../src/picorv32.v(1764)
  AL_MUX \picorv32_core/mux131_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/cpu_state [0]),
    .sel(\picorv32_core/mux131_b0_sel_is_1_o ),
    .o(\picorv32_core/n549 [0]));
  and \picorv32_core/mux131_b0_sel_is_1  (\picorv32_core/mux131_b0_sel_is_1_o , \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu , \picorv32_core/mem_done_neg );
  AL_MUX \picorv32_core/mux131_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/cpu_state [1]),
    .sel(\picorv32_core/mux131_b0_sel_is_1_o ),
    .o(\picorv32_core/n549 [1]));
  AL_MUX \picorv32_core/mux131_b2  (
    .i0(1'b0),
    .i1(\picorv32_core/cpu_state [2]),
    .sel(\picorv32_core/mux131_b0_sel_is_1_o ),
    .o(\picorv32_core/n549 [2]));
  AL_MUX \picorv32_core/mux131_b3  (
    .i0(1'b0),
    .i1(\picorv32_core/cpu_state [3]),
    .sel(\picorv32_core/mux131_b0_sel_is_1_o ),
    .o(\picorv32_core/n549 [3]));
  AL_MUX \picorv32_core/mux131_b4  (
    .i0(1'b0),
    .i1(\picorv32_core/cpu_state [4]),
    .sel(\picorv32_core/mux131_b0_sel_is_1_o ),
    .o(\picorv32_core/n549 [4]));
  AL_MUX \picorv32_core/mux131_b5  (
    .i0(1'b0),
    .i1(\picorv32_core/cpu_state [5]),
    .sel(\picorv32_core/mux131_b0_sel_is_1_o ),
    .o(\picorv32_core/n549 [5]));
  AL_MUX \picorv32_core/mux131_b6  (
    .i0(1'b1),
    .i1(\picorv32_core/cpu_state [6]),
    .sel(\picorv32_core/mux131_b0_sel_is_1_o ),
    .o(\picorv32_core/n549 [6]));
  AL_MUX \picorv32_core/mux131_b7  (
    .i0(1'b0),
    .i1(\picorv32_core/cpu_state [7]),
    .sel(\picorv32_core/mux131_b0_sel_is_1_o ),
    .o(\picorv32_core/n549 [7]));
  AL_MUX \picorv32_core/mux132_b0  (
    .i0(\picorv32_core/pcpi_rs1$0$ ),
    .i1(\picorv32_core/n576 [0]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [0]));
  and \picorv32_core/mux132_b0_sel_is_3  (\picorv32_core/mux132_b0_sel_is_3_o , \picorv32_core/n597 , \picorv32_core/n598 );
  AL_MUX \picorv32_core/mux132_b1  (
    .i0(\picorv32_core/pcpi_rs1$1$ ),
    .i1(\picorv32_core/n576 [1]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [1]));
  AL_MUX \picorv32_core/mux132_b10  (
    .i0(\picorv32_core/pcpi_rs1$10$ ),
    .i1(\picorv32_core/n576 [10]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [10]));
  AL_MUX \picorv32_core/mux132_b11  (
    .i0(\picorv32_core/pcpi_rs1$11$ ),
    .i1(\picorv32_core/n576 [11]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [11]));
  AL_MUX \picorv32_core/mux132_b12  (
    .i0(\picorv32_core/pcpi_rs1$12$ ),
    .i1(\picorv32_core/n576 [12]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [12]));
  AL_MUX \picorv32_core/mux132_b13  (
    .i0(\picorv32_core/pcpi_rs1$13$ ),
    .i1(\picorv32_core/n576 [13]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [13]));
  AL_MUX \picorv32_core/mux132_b14  (
    .i0(\picorv32_core/pcpi_rs1$14$ ),
    .i1(\picorv32_core/n576 [14]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [14]));
  AL_MUX \picorv32_core/mux132_b15  (
    .i0(\picorv32_core/pcpi_rs1$15$ ),
    .i1(\picorv32_core/n576 [15]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [15]));
  AL_MUX \picorv32_core/mux132_b16  (
    .i0(\picorv32_core/pcpi_rs1$16$ ),
    .i1(\picorv32_core/n576 [16]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [16]));
  AL_MUX \picorv32_core/mux132_b17  (
    .i0(\picorv32_core/pcpi_rs1$17$ ),
    .i1(\picorv32_core/n576 [17]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [17]));
  AL_MUX \picorv32_core/mux132_b18  (
    .i0(\picorv32_core/pcpi_rs1$18$ ),
    .i1(\picorv32_core/n576 [18]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [18]));
  AL_MUX \picorv32_core/mux132_b19  (
    .i0(\picorv32_core/pcpi_rs1$19$ ),
    .i1(\picorv32_core/n576 [19]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [19]));
  AL_MUX \picorv32_core/mux132_b2  (
    .i0(\picorv32_core/pcpi_rs1$2$ ),
    .i1(\picorv32_core/n576 [2]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [2]));
  AL_MUX \picorv32_core/mux132_b20  (
    .i0(\picorv32_core/pcpi_rs1$20$ ),
    .i1(\picorv32_core/n576 [20]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [20]));
  AL_MUX \picorv32_core/mux132_b21  (
    .i0(\picorv32_core/pcpi_rs1$21$ ),
    .i1(\picorv32_core/n576 [21]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [21]));
  AL_MUX \picorv32_core/mux132_b22  (
    .i0(\picorv32_core/pcpi_rs1$22$ ),
    .i1(\picorv32_core/n576 [22]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [22]));
  AL_MUX \picorv32_core/mux132_b23  (
    .i0(\picorv32_core/pcpi_rs1$23$ ),
    .i1(\picorv32_core/n576 [23]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [23]));
  AL_MUX \picorv32_core/mux132_b24  (
    .i0(\picorv32_core/pcpi_rs1$24$ ),
    .i1(\picorv32_core/n576 [24]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [24]));
  AL_MUX \picorv32_core/mux132_b25  (
    .i0(\picorv32_core/pcpi_rs1$25$ ),
    .i1(\picorv32_core/n576 [25]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [25]));
  AL_MUX \picorv32_core/mux132_b26  (
    .i0(\picorv32_core/pcpi_rs1$26$ ),
    .i1(\picorv32_core/n576 [26]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [26]));
  AL_MUX \picorv32_core/mux132_b27  (
    .i0(\picorv32_core/pcpi_rs1$27$ ),
    .i1(\picorv32_core/n576 [27]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [27]));
  AL_MUX \picorv32_core/mux132_b28  (
    .i0(\picorv32_core/pcpi_rs1$28$ ),
    .i1(\picorv32_core/n576 [28]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [28]));
  AL_MUX \picorv32_core/mux132_b29  (
    .i0(\picorv32_core/pcpi_rs1$29$ ),
    .i1(\picorv32_core/n576 [29]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [29]));
  AL_MUX \picorv32_core/mux132_b3  (
    .i0(\picorv32_core/pcpi_rs1$3$ ),
    .i1(\picorv32_core/n576 [3]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [3]));
  AL_MUX \picorv32_core/mux132_b30  (
    .i0(\picorv32_core/pcpi_rs1$30$ ),
    .i1(\picorv32_core/n576 [30]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [30]));
  AL_MUX \picorv32_core/mux132_b31  (
    .i0(\picorv32_core/pcpi_rs1$31$ ),
    .i1(\picorv32_core/n576 [31]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [31]));
  AL_MUX \picorv32_core/mux132_b32  (
    .i0(\picorv32_core/pcpi_rs1$0$ ),
    .i1(\picorv32_core/n576 [0]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [0]));
  and \picorv32_core/mux132_b32_sel_is_3  (\picorv32_core/mux132_b32_sel_is_3_o , \picorv32_core/n597 , \picorv32_core/n574 );
  AL_MUX \picorv32_core/mux132_b33  (
    .i0(\picorv32_core/pcpi_rs1$1$ ),
    .i1(\picorv32_core/n576 [1]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [1]));
  AL_MUX \picorv32_core/mux132_b34  (
    .i0(\picorv32_core/pcpi_rs1$2$ ),
    .i1(\picorv32_core/n576 [2]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [2]));
  AL_MUX \picorv32_core/mux132_b35  (
    .i0(\picorv32_core/pcpi_rs1$3$ ),
    .i1(\picorv32_core/n576 [3]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [3]));
  AL_MUX \picorv32_core/mux132_b36  (
    .i0(\picorv32_core/pcpi_rs1$4$ ),
    .i1(\picorv32_core/n576 [4]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [4]));
  AL_MUX \picorv32_core/mux132_b37  (
    .i0(\picorv32_core/pcpi_rs1$5$ ),
    .i1(\picorv32_core/n576 [5]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [5]));
  AL_MUX \picorv32_core/mux132_b38  (
    .i0(\picorv32_core/pcpi_rs1$6$ ),
    .i1(\picorv32_core/n576 [6]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [6]));
  AL_MUX \picorv32_core/mux132_b39  (
    .i0(\picorv32_core/pcpi_rs1$7$ ),
    .i1(\picorv32_core/n576 [7]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [7]));
  AL_MUX \picorv32_core/mux132_b4  (
    .i0(\picorv32_core/pcpi_rs1$4$ ),
    .i1(\picorv32_core/n576 [4]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [4]));
  AL_MUX \picorv32_core/mux132_b40  (
    .i0(\picorv32_core/pcpi_rs1$8$ ),
    .i1(\picorv32_core/n576 [8]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [8]));
  AL_MUX \picorv32_core/mux132_b41  (
    .i0(\picorv32_core/pcpi_rs1$9$ ),
    .i1(\picorv32_core/n576 [9]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [9]));
  AL_MUX \picorv32_core/mux132_b42  (
    .i0(\picorv32_core/pcpi_rs1$10$ ),
    .i1(\picorv32_core/n576 [10]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [10]));
  AL_MUX \picorv32_core/mux132_b43  (
    .i0(\picorv32_core/pcpi_rs1$11$ ),
    .i1(\picorv32_core/n576 [11]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [11]));
  AL_MUX \picorv32_core/mux132_b44  (
    .i0(\picorv32_core/pcpi_rs1$12$ ),
    .i1(\picorv32_core/n576 [12]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [12]));
  AL_MUX \picorv32_core/mux132_b45  (
    .i0(\picorv32_core/pcpi_rs1$13$ ),
    .i1(\picorv32_core/n576 [13]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [13]));
  AL_MUX \picorv32_core/mux132_b46  (
    .i0(\picorv32_core/pcpi_rs1$14$ ),
    .i1(\picorv32_core/n576 [14]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [14]));
  AL_MUX \picorv32_core/mux132_b47  (
    .i0(\picorv32_core/pcpi_rs1$15$ ),
    .i1(\picorv32_core/n576 [15]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [15]));
  AL_MUX \picorv32_core/mux132_b48  (
    .i0(\picorv32_core/pcpi_rs1$16$ ),
    .i1(\picorv32_core/n576 [16]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [16]));
  AL_MUX \picorv32_core/mux132_b49  (
    .i0(\picorv32_core/pcpi_rs1$17$ ),
    .i1(\picorv32_core/n576 [17]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [17]));
  AL_MUX \picorv32_core/mux132_b5  (
    .i0(\picorv32_core/pcpi_rs1$5$ ),
    .i1(\picorv32_core/n576 [5]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [5]));
  AL_MUX \picorv32_core/mux132_b50  (
    .i0(\picorv32_core/pcpi_rs1$18$ ),
    .i1(\picorv32_core/n576 [18]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [18]));
  AL_MUX \picorv32_core/mux132_b51  (
    .i0(\picorv32_core/pcpi_rs1$19$ ),
    .i1(\picorv32_core/n576 [19]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [19]));
  AL_MUX \picorv32_core/mux132_b52  (
    .i0(\picorv32_core/pcpi_rs1$20$ ),
    .i1(\picorv32_core/n576 [20]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [20]));
  AL_MUX \picorv32_core/mux132_b53  (
    .i0(\picorv32_core/pcpi_rs1$21$ ),
    .i1(\picorv32_core/n576 [21]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [21]));
  AL_MUX \picorv32_core/mux132_b54  (
    .i0(\picorv32_core/pcpi_rs1$22$ ),
    .i1(\picorv32_core/n576 [22]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [22]));
  AL_MUX \picorv32_core/mux132_b55  (
    .i0(\picorv32_core/pcpi_rs1$23$ ),
    .i1(\picorv32_core/n576 [23]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [23]));
  AL_MUX \picorv32_core/mux132_b56  (
    .i0(\picorv32_core/pcpi_rs1$24$ ),
    .i1(\picorv32_core/n576 [24]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [24]));
  AL_MUX \picorv32_core/mux132_b57  (
    .i0(\picorv32_core/pcpi_rs1$25$ ),
    .i1(\picorv32_core/n576 [25]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [25]));
  AL_MUX \picorv32_core/mux132_b58  (
    .i0(\picorv32_core/pcpi_rs1$26$ ),
    .i1(\picorv32_core/n576 [26]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [26]));
  AL_MUX \picorv32_core/mux132_b59  (
    .i0(\picorv32_core/pcpi_rs1$27$ ),
    .i1(\picorv32_core/n576 [27]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [27]));
  AL_MUX \picorv32_core/mux132_b6  (
    .i0(\picorv32_core/pcpi_rs1$6$ ),
    .i1(\picorv32_core/n576 [6]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [6]));
  AL_MUX \picorv32_core/mux132_b60  (
    .i0(\picorv32_core/pcpi_rs1$28$ ),
    .i1(\picorv32_core/n576 [28]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [28]));
  AL_MUX \picorv32_core/mux132_b61  (
    .i0(\picorv32_core/pcpi_rs1$29$ ),
    .i1(\picorv32_core/n576 [29]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [29]));
  AL_MUX \picorv32_core/mux132_b62  (
    .i0(\picorv32_core/pcpi_rs1$30$ ),
    .i1(\picorv32_core/n576 [30]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [30]));
  AL_MUX \picorv32_core/mux132_b63  (
    .i0(\picorv32_core/pcpi_rs1$31$ ),
    .i1(\picorv32_core/n576 [31]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n584 [31]));
  AL_MUX \picorv32_core/mux132_b7  (
    .i0(\picorv32_core/pcpi_rs1$7$ ),
    .i1(\picorv32_core/n576 [7]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [7]));
  AL_MUX \picorv32_core/mux132_b8  (
    .i0(\picorv32_core/pcpi_rs1$8$ ),
    .i1(\picorv32_core/n576 [8]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [8]));
  AL_MUX \picorv32_core/mux132_b9  (
    .i0(\picorv32_core/pcpi_rs1$9$ ),
    .i1(\picorv32_core/n576 [9]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n656 [9]));
  binary_mux_s1_w1 \picorv32_core/mux133_b0  (
    .i0(\picorv32_core/n563 [0]),
    .i1(\picorv32_core/n558 [0]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [0]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b1  (
    .i0(\picorv32_core/n563 [1]),
    .i1(\picorv32_core/n558 [1]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [1]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b10  (
    .i0(\picorv32_core/n563 [10]),
    .i1(\picorv32_core/n558 [10]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [10]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b11  (
    .i0(\picorv32_core/n563 [11]),
    .i1(\picorv32_core/n558 [11]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [11]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b12  (
    .i0(\picorv32_core/n563 [12]),
    .i1(\picorv32_core/n558 [12]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [12]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b13  (
    .i0(\picorv32_core/n563 [13]),
    .i1(\picorv32_core/n558 [13]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [13]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b14  (
    .i0(\picorv32_core/n563 [14]),
    .i1(\picorv32_core/n558 [14]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [14]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b15  (
    .i0(\picorv32_core/n563 [15]),
    .i1(\picorv32_core/n558 [15]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [15]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b16  (
    .i0(\picorv32_core/n563 [16]),
    .i1(\picorv32_core/n558 [16]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [16]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b17  (
    .i0(\picorv32_core/n563 [17]),
    .i1(\picorv32_core/n558 [17]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [17]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b18  (
    .i0(\picorv32_core/n563 [18]),
    .i1(\picorv32_core/n558 [18]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [18]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b19  (
    .i0(\picorv32_core/n563 [19]),
    .i1(\picorv32_core/n558 [19]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [19]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b2  (
    .i0(\picorv32_core/n563 [2]),
    .i1(\picorv32_core/n558 [2]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [2]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b20  (
    .i0(\picorv32_core/n563 [20]),
    .i1(\picorv32_core/n558 [20]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [20]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b21  (
    .i0(\picorv32_core/n563 [21]),
    .i1(\picorv32_core/n558 [21]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [21]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b22  (
    .i0(\picorv32_core/n563 [22]),
    .i1(\picorv32_core/n558 [22]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [22]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b23  (
    .i0(\picorv32_core/n563 [23]),
    .i1(\picorv32_core/n558 [23]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [23]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b24  (
    .i0(\picorv32_core/n563 [24]),
    .i1(\picorv32_core/n558 [24]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [24]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b25  (
    .i0(\picorv32_core/n563 [25]),
    .i1(\picorv32_core/n558 [25]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [25]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b26  (
    .i0(\picorv32_core/n563 [26]),
    .i1(\picorv32_core/n558 [26]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [26]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b27  (
    .i0(\picorv32_core/n563 [27]),
    .i1(\picorv32_core/n558 [27]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [27]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b28  (
    .i0(\picorv32_core/n563 [28]),
    .i1(\picorv32_core/n558 [28]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [28]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b29  (
    .i0(\picorv32_core/n563 [29]),
    .i1(\picorv32_core/n558 [29]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [29]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b3  (
    .i0(\picorv32_core/n563 [3]),
    .i1(\picorv32_core/n558 [3]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [3]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b30  (
    .i0(\picorv32_core/n563 [30]),
    .i1(\picorv32_core/n558 [30]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [30]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b31  (
    .i0(\picorv32_core/n563 [31]),
    .i1(\picorv32_core/n558 [31]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [31]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b4  (
    .i0(\picorv32_core/n563 [4]),
    .i1(\picorv32_core/n558 [4]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [4]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b5  (
    .i0(\picorv32_core/n563 [5]),
    .i1(\picorv32_core/n558 [5]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [5]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b6  (
    .i0(\picorv32_core/n563 [6]),
    .i1(\picorv32_core/n558 [6]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [6]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b7  (
    .i0(\picorv32_core/n563 [7]),
    .i1(\picorv32_core/n558 [7]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [7]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b8  (
    .i0(\picorv32_core/n563 [8]),
    .i1(\picorv32_core/n558 [8]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [8]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux133_b9  (
    .i0(\picorv32_core/n563 [9]),
    .i1(\picorv32_core/n558 [9]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n565 [9]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux134_b0  (
    .i0(\picorv32_core/n564 [0]),
    .i1(\picorv32_core/n559 [0]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n566 [0]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux134_b1  (
    .i0(\picorv32_core/n564 [1]),
    .i1(\picorv32_core/n559 [1]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n566 [1]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux134_b2  (
    .i0(\picorv32_core/n564 [2]),
    .i1(\picorv32_core/n559 [2]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n566 [2]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux134_b3  (
    .i0(\picorv32_core/n564 [3]),
    .i1(\picorv32_core/n559 [3]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n566 [3]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux134_b4  (
    .i0(\picorv32_core/n564 [4]),
    .i1(\picorv32_core/n559 [4]),
    .sel(\picorv32_core/n554 ),
    .o(\picorv32_core/n566 [4]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b0  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$0$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [0]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b1  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$1$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [1]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b10  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$10$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [10]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b11  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$11$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [11]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b12  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$12$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [12]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b13  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$13$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [13]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b14  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$14$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [14]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b15  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$15$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [15]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b16  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$16$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [16]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b17  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$17$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [17]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b18  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$18$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [18]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b19  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$19$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [19]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b2  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$2$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [2]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b20  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$20$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [20]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b21  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$21$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [21]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b22  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$22$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [22]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b23  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$23$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [23]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b24  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$24$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [24]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b25  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$25$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [25]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b26  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$26$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [26]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b27  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$27$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [27]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b28  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$28$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [28]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b29  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$29$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [29]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b3  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$3$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [3]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b30  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$30$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [30]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b31  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$31$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [31]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b4  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$4$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [4]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b5  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$5$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [5]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b6  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$6$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [6]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b7  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$7$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [7]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b8  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$8$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [8]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux135_b9  (
    .i0(1'bx),
    .i1(\picorv32_core/pcpi_rs1$9$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n567 [9]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux136_b0  (
    .i0(\picorv32_core/cpu_state [0]),
    .i1(1'b0),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n569 [0]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux136_b1  (
    .i0(\picorv32_core/cpu_state [1]),
    .i1(1'b0),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n569 [1]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux136_b2  (
    .i0(\picorv32_core/cpu_state [2]),
    .i1(1'b0),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n569 [2]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux136_b3  (
    .i0(\picorv32_core/cpu_state [3]),
    .i1(1'b0),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n569 [3]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux136_b4  (
    .i0(\picorv32_core/cpu_state [4]),
    .i1(1'b0),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n569 [4]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux136_b5  (
    .i0(\picorv32_core/cpu_state [5]),
    .i1(1'b0),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n569 [5]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux136_b6  (
    .i0(\picorv32_core/cpu_state [6]),
    .i1(1'b1),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n569 [6]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux136_b7  (
    .i0(\picorv32_core/cpu_state [7]),
    .i1(1'b0),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n569 [7]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b0  (
    .i0(\picorv32_core/n565 [0]),
    .i1(\picorv32_core/pcpi_rs1$0$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [0]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b1  (
    .i0(\picorv32_core/n565 [1]),
    .i1(\picorv32_core/pcpi_rs1$1$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [1]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b10  (
    .i0(\picorv32_core/n565 [10]),
    .i1(\picorv32_core/pcpi_rs1$10$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [10]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b11  (
    .i0(\picorv32_core/n565 [11]),
    .i1(\picorv32_core/pcpi_rs1$11$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [11]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b12  (
    .i0(\picorv32_core/n565 [12]),
    .i1(\picorv32_core/pcpi_rs1$12$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [12]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b13  (
    .i0(\picorv32_core/n565 [13]),
    .i1(\picorv32_core/pcpi_rs1$13$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [13]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b14  (
    .i0(\picorv32_core/n565 [14]),
    .i1(\picorv32_core/pcpi_rs1$14$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [14]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b15  (
    .i0(\picorv32_core/n565 [15]),
    .i1(\picorv32_core/pcpi_rs1$15$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [15]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b16  (
    .i0(\picorv32_core/n565 [16]),
    .i1(\picorv32_core/pcpi_rs1$16$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [16]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b17  (
    .i0(\picorv32_core/n565 [17]),
    .i1(\picorv32_core/pcpi_rs1$17$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [17]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b18  (
    .i0(\picorv32_core/n565 [18]),
    .i1(\picorv32_core/pcpi_rs1$18$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [18]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b19  (
    .i0(\picorv32_core/n565 [19]),
    .i1(\picorv32_core/pcpi_rs1$19$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [19]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b2  (
    .i0(\picorv32_core/n565 [2]),
    .i1(\picorv32_core/pcpi_rs1$2$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [2]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b20  (
    .i0(\picorv32_core/n565 [20]),
    .i1(\picorv32_core/pcpi_rs1$20$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [20]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b21  (
    .i0(\picorv32_core/n565 [21]),
    .i1(\picorv32_core/pcpi_rs1$21$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [21]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b22  (
    .i0(\picorv32_core/n565 [22]),
    .i1(\picorv32_core/pcpi_rs1$22$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [22]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b23  (
    .i0(\picorv32_core/n565 [23]),
    .i1(\picorv32_core/pcpi_rs1$23$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [23]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b24  (
    .i0(\picorv32_core/n565 [24]),
    .i1(\picorv32_core/pcpi_rs1$24$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [24]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b25  (
    .i0(\picorv32_core/n565 [25]),
    .i1(\picorv32_core/pcpi_rs1$25$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [25]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b26  (
    .i0(\picorv32_core/n565 [26]),
    .i1(\picorv32_core/pcpi_rs1$26$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [26]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b27  (
    .i0(\picorv32_core/n565 [27]),
    .i1(\picorv32_core/pcpi_rs1$27$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [27]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b28  (
    .i0(\picorv32_core/n565 [28]),
    .i1(\picorv32_core/pcpi_rs1$28$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [28]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b29  (
    .i0(\picorv32_core/n565 [29]),
    .i1(\picorv32_core/pcpi_rs1$29$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [29]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b3  (
    .i0(\picorv32_core/n565 [3]),
    .i1(\picorv32_core/pcpi_rs1$3$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [3]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b30  (
    .i0(\picorv32_core/n565 [30]),
    .i1(\picorv32_core/pcpi_rs1$30$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [30]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b31  (
    .i0(\picorv32_core/n565 [31]),
    .i1(\picorv32_core/pcpi_rs1$31$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [31]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b4  (
    .i0(\picorv32_core/n565 [4]),
    .i1(\picorv32_core/pcpi_rs1$4$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [4]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b5  (
    .i0(\picorv32_core/n565 [5]),
    .i1(\picorv32_core/pcpi_rs1$5$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [5]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b6  (
    .i0(\picorv32_core/n565 [6]),
    .i1(\picorv32_core/pcpi_rs1$6$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [6]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b7  (
    .i0(\picorv32_core/n565 [7]),
    .i1(\picorv32_core/pcpi_rs1$7$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [7]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b8  (
    .i0(\picorv32_core/n565 [8]),
    .i1(\picorv32_core/pcpi_rs1$8$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [8]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux137_b9  (
    .i0(\picorv32_core/n565 [9]),
    .i1(\picorv32_core/pcpi_rs1$9$ ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n570 [9]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux138_b0  (
    .i0(\picorv32_core/n566 [0]),
    .i1(1'bx),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n571 [0]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux138_b1  (
    .i0(\picorv32_core/n566 [1]),
    .i1(1'bx),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n571 [1]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux138_b2  (
    .i0(\picorv32_core/n566 [2]),
    .i1(1'bx),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n571 [2]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux138_b3  (
    .i0(\picorv32_core/n566 [3]),
    .i1(1'bx),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n571 [3]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux138_b4  (
    .i0(\picorv32_core/n566 [4]),
    .i1(1'bx),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n571 [4]));  // ../src/picorv32.v(1789)
  binary_mux_s1_w1 \picorv32_core/mux13_b0  (
    .i0(\picorv32_core/n66 [0]),
    .i1(1'b1),
    .sel(\picorv32_core/n67 ),
    .o(\picorv32_core/n68 [0]));  // ../src/picorv32.v(454)
  AL_MUX \picorv32_core/mux13_b1  (
    .i0(1'b1),
    .i1(\picorv32_core/n64 [1]),
    .sel(\picorv32_core/mux13_b1_sel_is_0_o ),
    .o(\picorv32_core/n68 [1]));
  and \picorv32_core/mux13_b1_sel_is_0  (\picorv32_core/mux13_b1_sel_is_0_o , \picorv32_core/n67_neg , \picorv32_core/n65_neg );
  AL_MUX \picorv32_core/mux13_b2  (
    .i0(1'b1),
    .i1(\picorv32_core/n62 [2]),
    .sel(\picorv32_core/mux13_b2_sel_is_2_o ),
    .o(\picorv32_core/n68 [2]));
  and \picorv32_core/mux13_b2_sel_is_2  (\picorv32_core/mux13_b2_sel_is_2_o , \picorv32_core/n67_neg , \picorv32_core/mux20_b2_sel_is_0_o );
  binary_mux_s1_w1 \picorv32_core/mux142_b0  (
    .i0(\picorv32_core/n42 [7]),
    .i1(1'b0),
    .sel(\picorv32_core/n99 ),
    .o(\picorv32_core/n52 [0]));  // ../src/picorv32.v(504)
  binary_mux_s1_w1 \picorv32_core/mux142_b1  (
    .i0(\picorv32_core/n42 [8]),
    .i1(1'b0),
    .sel(\picorv32_core/n99 ),
    .o(\picorv32_core/n52 [1]));  // ../src/picorv32.v(504)
  binary_mux_s1_w1 \picorv32_core/mux142_b2  (
    .i0(\picorv32_core/n42 [9]),
    .i1(\picorv32_core/mem_rdata_latched [6]),
    .sel(\picorv32_core/n99 ),
    .o(\picorv32_core/n52 [2]));  // ../src/picorv32.v(504)
  binary_mux_s1_w1 \picorv32_core/mux142_b3  (
    .i0(\picorv32_core/n42 [10]),
    .i1(\picorv32_core/mem_rdata_latched [10]),
    .sel(\picorv32_core/n99 ),
    .o(\picorv32_core/n52 [3]));  // ../src/picorv32.v(504)
  binary_mux_s1_w1 \picorv32_core/mux142_b4  (
    .i0(\picorv32_core/n42 [11]),
    .i1(\picorv32_core/mem_rdata_latched [11]),
    .sel(\picorv32_core/n99 ),
    .o(\picorv32_core/n52 [4]));  // ../src/picorv32.v(504)
  binary_mux_s1_w1 \picorv32_core/mux142_b7  (
    .i0(\picorv32_core/n42 [9]),
    .i1(\picorv32_core/mem_rdata_latched [9]),
    .sel(\picorv32_core/n99 ),
    .o(\picorv32_core/n108 [2]));  // ../src/picorv32.v(504)
  AL_MUX \picorv32_core/mux143_b0  (
    .i0(\picorv32_core/mem_wordsize [0]),
    .i1(\picorv32_core/n601 [0]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n652 [0]));
  AL_MUX \picorv32_core/mux143_b1  (
    .i0(\picorv32_core/mem_wordsize [1]),
    .i1(\picorv32_core/n601 [1]),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n652 [1]));
  AL_MUX \picorv32_core/mux143_b2  (
    .i0(\picorv32_core/mem_wordsize [0]),
    .i1(\picorv32_core/n575 [0]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n583 [0]));
  AL_MUX \picorv32_core/mux143_b3  (
    .i0(\picorv32_core/mem_wordsize [1]),
    .i1(\picorv32_core/n575 [1]),
    .sel(\picorv32_core/mux132_b32_sel_is_3_o ),
    .o(\picorv32_core/n583 [1]));
  binary_mux_s1_w1 \picorv32_core/mux146_b0  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [0]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [0]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b1  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [1]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [1]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b10  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [10]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [10]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b11  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [11]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [11]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b12  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [12]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [12]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b13  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [13]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [13]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b14  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [14]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [14]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b15  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [15]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [15]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b16  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [16]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [16]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b17  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [17]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [17]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b18  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [18]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [18]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b19  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [19]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [19]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b2  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [2]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [2]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b20  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [20]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [20]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b21  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [21]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [21]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b22  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [22]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [22]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b23  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [23]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [23]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b24  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [24]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [24]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b25  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [25]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [25]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b26  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [26]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [26]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b27  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [27]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [27]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b28  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [28]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [28]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b29  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [29]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [29]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b3  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [3]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [3]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b30  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [30]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [30]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b31  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [31]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [31]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b4  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [4]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [4]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b5  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [5]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [5]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b6  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [6]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [6]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b7  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [7]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [7]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b8  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [8]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [8]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux146_b9  (
    .i0(1'bx),
    .i1(\picorv32_core/n641 [9]),
    .sel(\picorv32_core/n580 ),
    .o(\picorv32_core/n642 [9]));  // ../src/picorv32.v(1848)
  binary_mux_s1_w1 \picorv32_core/mux147_b0  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [0]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [0]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b1  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [1]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [1]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b10  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [10]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [10]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b11  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [11]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [11]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b12  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [12]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [12]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b13  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [13]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [13]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b14  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [14]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [14]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b15  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [15]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [15]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b16  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [16]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [16]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b17  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [17]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [17]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b18  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [18]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [18]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b19  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [19]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [19]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b2  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [2]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [2]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b20  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [20]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [20]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b21  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [21]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [21]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b22  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [22]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [22]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b23  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [23]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [23]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b24  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [24]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [24]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b25  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [25]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [25]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b26  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [26]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [26]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b27  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [27]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [27]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b28  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [28]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [28]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b29  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [29]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [29]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b3  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [3]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [3]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b30  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [30]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [30]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b31  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [31]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [31]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b4  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [4]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [4]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b5  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [5]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [5]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b6  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [6]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [6]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b7  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [7]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [7]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b8  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [8]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [8]));  // ../src/picorv32.v(1849)
  binary_mux_s1_w1 \picorv32_core/mux147_b9  (
    .i0(1'bx),
    .i1(\picorv32_core/n642 [9]),
    .sel(\picorv32_core/n597 ),
    .o(\picorv32_core/n658 [9]));  // ../src/picorv32.v(1849)
  AL_MUX \picorv32_core/mux148_b0  (
    .i0(\picorv32_core/cpu_state [0]),
    .i1(1'b0),
    .sel(\picorv32_core/mux148_b0_sel_is_3_o ),
    .o(\picorv32_core/n661 [0]));
  and \picorv32_core/mux148_b0_sel_is_3  (\picorv32_core/mux148_b0_sel_is_3_o , \picorv32_core/n597 , \picorv32_core/n580 );
  AL_MUX \picorv32_core/mux148_b1  (
    .i0(\picorv32_core/cpu_state [1]),
    .i1(1'b0),
    .sel(\picorv32_core/mux148_b0_sel_is_3_o ),
    .o(\picorv32_core/n661 [1]));
  AL_MUX \picorv32_core/mux148_b2  (
    .i0(\picorv32_core/cpu_state [2]),
    .i1(1'b0),
    .sel(\picorv32_core/mux148_b0_sel_is_3_o ),
    .o(\picorv32_core/n661 [2]));
  AL_MUX \picorv32_core/mux148_b3  (
    .i0(\picorv32_core/cpu_state [3]),
    .i1(1'b0),
    .sel(\picorv32_core/mux148_b0_sel_is_3_o ),
    .o(\picorv32_core/n661 [3]));
  AL_MUX \picorv32_core/mux148_b4  (
    .i0(\picorv32_core/cpu_state [4]),
    .i1(1'b0),
    .sel(\picorv32_core/mux148_b0_sel_is_3_o ),
    .o(\picorv32_core/n661 [4]));
  AL_MUX \picorv32_core/mux148_b5  (
    .i0(\picorv32_core/cpu_state [5]),
    .i1(1'b0),
    .sel(\picorv32_core/mux148_b0_sel_is_3_o ),
    .o(\picorv32_core/n661 [5]));
  AL_MUX \picorv32_core/mux148_b6  (
    .i0(\picorv32_core/cpu_state [6]),
    .i1(1'b1),
    .sel(\picorv32_core/mux148_b0_sel_is_3_o ),
    .o(\picorv32_core/n661 [6]));
  AL_MUX \picorv32_core/mux148_b7  (
    .i0(\picorv32_core/cpu_state [7]),
    .i1(1'b0),
    .sel(\picorv32_core/mux148_b0_sel_is_3_o ),
    .o(\picorv32_core/n661 [7]));
  binary_mux_s1_w1 \picorv32_core/mux14_b8  (
    .i0(\picorv32_core/n42 [30]),
    .i1(1'b0),
    .sel(\picorv32_core/n54 ),
    .o(\picorv32_core/n55 [8]));  // ../src/picorv32.v(441)
  binary_mux_s1_w1 \picorv32_core/mux154_b0  (
    .i0(\picorv32_core/n692 [0]),
    .i1(1'b0),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n716 [0]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux154_b1  (
    .i0(\picorv32_core/n692 [1]),
    .i1(1'b0),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n716 [1]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux154_b2  (
    .i0(\picorv32_core/n692 [2]),
    .i1(1'b0),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n716 [2]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux154_b3  (
    .i0(\picorv32_core/n692 [3]),
    .i1(1'b0),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n716 [3]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux154_b4  (
    .i0(\picorv32_core/n692 [4]),
    .i1(1'b0),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n716 [4]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux154_b5  (
    .i0(\picorv32_core/n692 [5]),
    .i1(1'b0),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n716 [5]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux154_b7  (
    .i0(\picorv32_core/n692 [7]),
    .i1(1'b0),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n716 [7]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b0  (
    .i0(\picorv32_core/n695 [0]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [0]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b1  (
    .i0(\picorv32_core/n695 [1]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [1]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b10  (
    .i0(\picorv32_core/n695 [10]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [10]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b11  (
    .i0(\picorv32_core/n695 [11]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [11]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b12  (
    .i0(\picorv32_core/n695 [12]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [12]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b13  (
    .i0(\picorv32_core/n695 [13]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [13]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b14  (
    .i0(\picorv32_core/n695 [14]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [14]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b15  (
    .i0(\picorv32_core/n695 [15]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [15]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b16  (
    .i0(\picorv32_core/n695 [16]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [16]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b17  (
    .i0(\picorv32_core/n695 [17]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [17]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b18  (
    .i0(\picorv32_core/n695 [18]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [18]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b19  (
    .i0(\picorv32_core/n695 [19]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [19]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b2  (
    .i0(\picorv32_core/n695 [2]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [2]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b20  (
    .i0(\picorv32_core/n695 [20]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [20]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b21  (
    .i0(\picorv32_core/n695 [21]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [21]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b22  (
    .i0(\picorv32_core/n695 [22]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [22]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b23  (
    .i0(\picorv32_core/n695 [23]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [23]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b24  (
    .i0(\picorv32_core/n695 [24]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [24]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b25  (
    .i0(\picorv32_core/n695 [25]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [25]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b26  (
    .i0(\picorv32_core/n695 [26]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [26]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b27  (
    .i0(\picorv32_core/n695 [27]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [27]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b28  (
    .i0(\picorv32_core/n695 [28]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [28]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b29  (
    .i0(\picorv32_core/n695 [29]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [29]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b3  (
    .i0(\picorv32_core/n695 [3]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [3]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b30  (
    .i0(\picorv32_core/n695 [30]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [30]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b31  (
    .i0(\picorv32_core/n695 [31]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [31]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b4  (
    .i0(\picorv32_core/n695 [4]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [4]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b5  (
    .i0(\picorv32_core/n695 [5]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [5]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b6  (
    .i0(\picorv32_core/n695 [6]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [6]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b7  (
    .i0(\picorv32_core/n695 [7]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [7]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b8  (
    .i0(\picorv32_core/n695 [8]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [8]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux159_b9  (
    .i0(\picorv32_core/n695 [9]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n725 [9]));  // ../src/picorv32.v(1851)
  and \picorv32_core/mux15_b0_sel_is_0  (\picorv32_core/mux15_b0_sel_is_0_o , \picorv32_core/n56_neg , \picorv32_core/n54_neg );
  AL_MUX \picorv32_core/mux15_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [13]),
    .sel(\picorv32_core/mux15_b0_sel_is_0_o ),
    .o(\picorv32_core/n57 [1]));
  AL_MUX \picorv32_core/mux15_b3  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [25]),
    .sel(\picorv32_core/mux15_b0_sel_is_0_o ),
    .o(\picorv32_core/n57 [3]));
  AL_MUX \picorv32_core/mux15_b4  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [26]),
    .sel(\picorv32_core/mux15_b0_sel_is_0_o ),
    .o(\picorv32_core/n57 [4]));
  AL_MUX \picorv32_core/mux15_b5  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [27]),
    .sel(\picorv32_core/mux15_b0_sel_is_0_o ),
    .o(\picorv32_core/n57 [5]));
  AL_MUX \picorv32_core/mux15_b6  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [28]),
    .sel(\picorv32_core/mux15_b0_sel_is_0_o ),
    .o(\picorv32_core/n57 [6]));
  AL_MUX \picorv32_core/mux15_b7  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [29]),
    .sel(\picorv32_core/mux15_b0_sel_is_0_o ),
    .o(\picorv32_core/n57 [7]));
  binary_mux_s1_w1 \picorv32_core/mux15_b8  (
    .i0(\picorv32_core/n55 [8]),
    .i1(1'b1),
    .sel(\picorv32_core/n56 ),
    .o(\picorv32_core/n57 [8]));  // ../src/picorv32.v(445)
  AL_MUX \picorv32_core/mux15_b9  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [31]),
    .sel(\picorv32_core/mux15_b0_sel_is_0_o ),
    .o(\picorv32_core/n57 [9]));
  binary_mux_s1_w1 \picorv32_core/mux160_b0  (
    .i0(\picorv32_core/n696 [0]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n726 [0]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux160_b1  (
    .i0(\picorv32_core/n696 [1]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n726 [1]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux160_b2  (
    .i0(\picorv32_core/n696 [2]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n726 [2]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux160_b3  (
    .i0(\picorv32_core/n696 [3]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n726 [3]));  // ../src/picorv32.v(1851)
  binary_mux_s1_w1 \picorv32_core/mux160_b4  (
    .i0(\picorv32_core/n696 [4]),
    .i1(1'bx),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n726 [4]));  // ../src/picorv32.v(1851)
  and \picorv32_core/mux162_b0_sel_is_0  (\picorv32_core/mux162_b0_sel_is_0_o , \picorv32_core/n740_neg , \picorv32_core/n736_neg );
  not \picorv32_core/mux162_b0_sel_is_0_o_inv  (\picorv32_core/mux162_b0_sel_is_0_o_neg , \picorv32_core/mux162_b0_sel_is_0_o );
  and \picorv32_core/mux163_b0_sel_is_1  (\picorv32_core/mux163_b0_sel_is_1_o , \picorv32_core/n733 , \picorv32_core/mux162_b0_sel_is_0_o_neg );
  not \picorv32_core/mux163_b0_sel_is_1_o_inv  (\picorv32_core/mux163_b0_sel_is_1_o_neg , \picorv32_core/mux163_b0_sel_is_1_o );
  and \picorv32_core/mux164_b0_sel_is_0  (\picorv32_core/mux164_b0_sel_is_0_o , \picorv32_core/n744_neg , \picorv32_core/mux163_b0_sel_is_1_o_neg );
  AL_MUX \picorv32_core/mux165_b0  (
    .i0(mem_la_wdata[0]),
    .i1(\picorv32_core/pcpi_rs2$16$ ),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(mem_la_wdata[16]));
  and \picorv32_core/mux165_b0_sel_is_0  (\picorv32_core/mux165_b0_sel_is_0_o , \picorv32_core/mem_wordsize$0$_neg , \picorv32_core/mem_wordsize$1$_neg );
  AL_MUX \picorv32_core/mux165_b1  (
    .i0(mem_la_wdata[1]),
    .i1(\picorv32_core/pcpi_rs2$17$ ),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(mem_la_wdata[17]));
  binary_mux_s2_w1 \picorv32_core/mux165_b10  (
    .i0(\picorv32_core/pcpi_rs2$26$ ),
    .i1(\picorv32_core/pcpi_rs2$10$ ),
    .i2(mem_la_wdata[2]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(mem_la_wdata[26]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux165_b11  (
    .i0(\picorv32_core/pcpi_rs2$27$ ),
    .i1(\picorv32_core/pcpi_rs2$11$ ),
    .i2(mem_la_wdata[3]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(mem_la_wdata[27]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux165_b12  (
    .i0(\picorv32_core/pcpi_rs2$28$ ),
    .i1(\picorv32_core/pcpi_rs2$12$ ),
    .i2(mem_la_wdata[4]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(mem_la_wdata[28]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux165_b13  (
    .i0(\picorv32_core/pcpi_rs2$29$ ),
    .i1(\picorv32_core/pcpi_rs2$13$ ),
    .i2(mem_la_wdata[5]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(mem_la_wdata[29]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux165_b14  (
    .i0(\picorv32_core/pcpi_rs2$30$ ),
    .i1(\picorv32_core/pcpi_rs2$14$ ),
    .i2(mem_la_wdata[6]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(mem_la_wdata[30]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux165_b15  (
    .i0(\picorv32_core/pcpi_rs2$31$ ),
    .i1(\picorv32_core/pcpi_rs2$15$ ),
    .i2(mem_la_wdata[7]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(mem_la_wdata[31]));  // ../src/picorv32.v(391)
  AL_MUX \picorv32_core/mux165_b2  (
    .i0(mem_la_wdata[2]),
    .i1(\picorv32_core/pcpi_rs2$18$ ),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(mem_la_wdata[18]));
  AL_MUX \picorv32_core/mux165_b3  (
    .i0(mem_la_wdata[3]),
    .i1(\picorv32_core/pcpi_rs2$19$ ),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(mem_la_wdata[19]));
  AL_MUX \picorv32_core/mux165_b4  (
    .i0(mem_la_wdata[4]),
    .i1(\picorv32_core/pcpi_rs2$20$ ),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(mem_la_wdata[20]));
  AL_MUX \picorv32_core/mux165_b5  (
    .i0(mem_la_wdata[5]),
    .i1(\picorv32_core/pcpi_rs2$21$ ),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(mem_la_wdata[21]));
  AL_MUX \picorv32_core/mux165_b6  (
    .i0(mem_la_wdata[6]),
    .i1(\picorv32_core/pcpi_rs2$22$ ),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(mem_la_wdata[22]));
  AL_MUX \picorv32_core/mux165_b7  (
    .i0(mem_la_wdata[7]),
    .i1(\picorv32_core/pcpi_rs2$23$ ),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(mem_la_wdata[23]));
  binary_mux_s2_w1 \picorv32_core/mux165_b8  (
    .i0(\picorv32_core/pcpi_rs2$24$ ),
    .i1(\picorv32_core/pcpi_rs2$8$ ),
    .i2(mem_la_wdata[0]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(mem_la_wdata[24]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux165_b9  (
    .i0(\picorv32_core/pcpi_rs2$25$ ),
    .i1(\picorv32_core/pcpi_rs2$9$ ),
    .i2(mem_la_wdata[1]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(mem_la_wdata[25]));  // ../src/picorv32.v(391)
  binary_mux_s1_w1 \picorv32_core/mux16_b0  (
    .i0(\picorv32_core/mem_rdata_latched [2]),
    .i1(1'b0),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n53 [0]));  // ../src/picorv32.v(435)
  binary_mux_s1_w1 \picorv32_core/mux16_b1  (
    .i0(\picorv32_core/mem_rdata_latched [3]),
    .i1(1'b0),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n53 [1]));  // ../src/picorv32.v(435)
  binary_mux_s1_w1 \picorv32_core/mux16_b10  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(1'b0),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n53 [10]));  // ../src/picorv32.v(435)
  binary_mux_s1_w1 \picorv32_core/mux16_b12  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/mem_rdata_latched [6]),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n53 [12]));  // ../src/picorv32.v(435)
  binary_mux_s1_w1 \picorv32_core/mux16_b13  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/mem_rdata_latched [2]),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n53 [13]));  // ../src/picorv32.v(435)
  binary_mux_s1_w1 \picorv32_core/mux16_b14  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/mem_rdata_latched [5]),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n53 [14]));  // ../src/picorv32.v(435)
  binary_mux_s1_w1 \picorv32_core/mux16_b15  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/mem_rdata_latched [3]),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n53 [15]));  // ../src/picorv32.v(435)
  binary_mux_s1_w1 \picorv32_core/mux16_b16  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/mem_rdata_latched [4]),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n53 [16]));  // ../src/picorv32.v(435)
  binary_mux_s1_w1 \picorv32_core/mux16_b2  (
    .i0(\picorv32_core/mem_rdata_latched [4]),
    .i1(1'b0),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n53 [2]));  // ../src/picorv32.v(435)
  binary_mux_s1_w1 \picorv32_core/mux17_b0  (
    .i0(\picorv32_core/n42 [20]),
    .i1(\picorv32_core/mem_rdata_latched [2]),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n60 [0]));  // ../src/picorv32.v(449)
  binary_mux_s1_w1 \picorv32_core/mux17_b1  (
    .i0(\picorv32_core/n42 [21]),
    .i1(\picorv32_core/mem_rdata_latched [3]),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n60 [1]));  // ../src/picorv32.v(449)
  binary_mux_s1_w1 \picorv32_core/mux17_b2  (
    .i0(\picorv32_core/n42 [22]),
    .i1(\picorv32_core/mem_rdata_latched [4]),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n60 [2]));  // ../src/picorv32.v(449)
  binary_mux_s1_w1 \picorv32_core/mux17_b3  (
    .i0(\picorv32_core/n42 [23]),
    .i1(\picorv32_core/mem_rdata_latched [5]),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n60 [3]));  // ../src/picorv32.v(449)
  binary_mux_s1_w1 \picorv32_core/mux17_b4  (
    .i0(\picorv32_core/n42 [24]),
    .i1(\picorv32_core/mem_rdata_latched [6]),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n60 [4]));  // ../src/picorv32.v(449)
  binary_mux_s1_w1 \picorv32_core/mux18_b2  (
    .i0(\picorv32_core/n59 [2]),
    .i1(1'b0),
    .sel(\picorv32_core/n61 ),
    .o(\picorv32_core/n62 [2]));  // ../src/picorv32.v(451)
  and \picorv32_core/mux19_b0_sel_is_0  (\picorv32_core/mux19_b0_sel_is_0_o , \picorv32_core/n63_neg , \picorv32_core/n61_neg );
  AL_MUX \picorv32_core/mux19_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/n59 [1]),
    .sel(\picorv32_core/mux19_b0_sel_is_0_o ),
    .o(\picorv32_core/n64 [1]));
  binary_mux_s1_w1 \picorv32_core/mux1_b0  (
    .i0(\picorv32_core/mem_rdata_q [0]),
    .i1(mem_rdata[0]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [0]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b1  (
    .i0(\picorv32_core/mem_rdata_q [1]),
    .i1(mem_rdata[1]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [1]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b10  (
    .i0(\picorv32_core/mem_rdata_q [10]),
    .i1(mem_rdata[10]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [10]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b11  (
    .i0(\picorv32_core/mem_rdata_q [11]),
    .i1(mem_rdata[11]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [11]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b12  (
    .i0(\picorv32_core/mem_rdata_q [12]),
    .i1(mem_rdata[12]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [12]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b13  (
    .i0(\picorv32_core/mem_rdata_q [13]),
    .i1(mem_rdata[13]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [13]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b14  (
    .i0(\picorv32_core/mem_rdata_q [14]),
    .i1(mem_rdata[14]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [14]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b15  (
    .i0(\picorv32_core/mem_rdata_q [15]),
    .i1(mem_rdata[15]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [15]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b16  (
    .i0(\picorv32_core/mem_rdata_q [16]),
    .i1(mem_rdata[16]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [16]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b17  (
    .i0(\picorv32_core/mem_rdata_q [17]),
    .i1(mem_rdata[17]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [17]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b18  (
    .i0(\picorv32_core/mem_rdata_q [18]),
    .i1(mem_rdata[18]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [18]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b19  (
    .i0(\picorv32_core/mem_rdata_q [19]),
    .i1(mem_rdata[19]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [19]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b2  (
    .i0(\picorv32_core/mem_rdata_q [2]),
    .i1(mem_rdata[2]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [2]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b20  (
    .i0(\picorv32_core/mem_rdata_q [20]),
    .i1(mem_rdata[20]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [20]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b21  (
    .i0(\picorv32_core/mem_rdata_q [21]),
    .i1(mem_rdata[21]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [21]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b22  (
    .i0(\picorv32_core/mem_rdata_q [22]),
    .i1(mem_rdata[22]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [22]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b23  (
    .i0(\picorv32_core/mem_rdata_q [23]),
    .i1(mem_rdata[23]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [23]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b24  (
    .i0(\picorv32_core/mem_rdata_q [24]),
    .i1(mem_rdata[24]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [24]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b25  (
    .i0(\picorv32_core/mem_rdata_q [25]),
    .i1(mem_rdata[25]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [25]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b26  (
    .i0(\picorv32_core/mem_rdata_q [26]),
    .i1(mem_rdata[26]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [26]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b27  (
    .i0(\picorv32_core/mem_rdata_q [27]),
    .i1(mem_rdata[27]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [27]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b28  (
    .i0(\picorv32_core/mem_rdata_q [28]),
    .i1(mem_rdata[28]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [28]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b29  (
    .i0(\picorv32_core/mem_rdata_q [29]),
    .i1(mem_rdata[29]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [29]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b3  (
    .i0(\picorv32_core/mem_rdata_q [3]),
    .i1(mem_rdata[3]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [3]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b30  (
    .i0(\picorv32_core/mem_rdata_q [30]),
    .i1(mem_rdata[30]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [30]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b31  (
    .i0(\picorv32_core/mem_rdata_q [31]),
    .i1(mem_rdata[31]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [31]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b4  (
    .i0(\picorv32_core/mem_rdata_q [4]),
    .i1(mem_rdata[4]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [4]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b5  (
    .i0(\picorv32_core/mem_rdata_q [5]),
    .i1(mem_rdata[5]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [5]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b6  (
    .i0(\picorv32_core/mem_rdata_q [6]),
    .i1(mem_rdata[6]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [6]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b7  (
    .i0(\picorv32_core/mem_rdata_q [7]),
    .i1(mem_rdata[7]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [7]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b8  (
    .i0(\picorv32_core/mem_rdata_q [8]),
    .i1(mem_rdata[8]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [8]));  // ../src/picorv32.v(348)
  binary_mux_s1_w1 \picorv32_core/mux1_b9  (
    .i0(\picorv32_core/mem_rdata_q [9]),
    .i1(mem_rdata[9]),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/mem_rdata_latched_noshuffle [9]));  // ../src/picorv32.v(348)
  AL_MUX \picorv32_core/mux20_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/n59 [0]),
    .sel(\picorv32_core/mux20_b0_sel_is_2_o ),
    .o(\picorv32_core/n66 [0]));
  and \picorv32_core/mux20_b0_sel_is_2  (\picorv32_core/mux20_b0_sel_is_2_o , \picorv32_core/n65_neg , \picorv32_core/mux19_b0_sel_is_0_o );
  and \picorv32_core/mux20_b2_sel_is_0  (\picorv32_core/mux20_b2_sel_is_0_o , \picorv32_core/n65_neg , \picorv32_core/n63_neg );
  AL_MUX \picorv32_core/mux21_b0  (
    .i0(1'b1),
    .i1(\picorv32_core/n42 [12]),
    .sel(\picorv32_core/mux21_b0_sel_is_2_o ),
    .o(\picorv32_core/n59 [0]));
  and \picorv32_core/mux21_b0_sel_is_2  (\picorv32_core/mux21_b0_sel_is_2_o , \picorv32_core/n58_neg , \picorv32_core/mux15_b0_sel_is_0_o );
  binary_mux_s1_w1 \picorv32_core/mux21_b1  (
    .i0(\picorv32_core/n57 [1]),
    .i1(1'b1),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n59 [1]));  // ../src/picorv32.v(449)
  AL_MUX \picorv32_core/mux21_b2  (
    .i0(1'b1),
    .i1(\picorv32_core/n42 [14]),
    .sel(\picorv32_core/mux21_b0_sel_is_2_o ),
    .o(\picorv32_core/n59 [2]));
  binary_mux_s1_w1 \picorv32_core/mux21_b3  (
    .i0(\picorv32_core/n57 [3]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n59 [3]));  // ../src/picorv32.v(449)
  binary_mux_s1_w1 \picorv32_core/mux21_b4  (
    .i0(\picorv32_core/n57 [4]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n59 [4]));  // ../src/picorv32.v(449)
  binary_mux_s1_w1 \picorv32_core/mux21_b5  (
    .i0(\picorv32_core/n57 [5]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n59 [5]));  // ../src/picorv32.v(449)
  binary_mux_s1_w1 \picorv32_core/mux21_b6  (
    .i0(\picorv32_core/n57 [6]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n59 [6]));  // ../src/picorv32.v(449)
  binary_mux_s1_w1 \picorv32_core/mux21_b7  (
    .i0(\picorv32_core/n57 [7]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n59 [7]));  // ../src/picorv32.v(449)
  binary_mux_s1_w1 \picorv32_core/mux21_b8  (
    .i0(\picorv32_core/n57 [8]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n59 [8]));  // ../src/picorv32.v(449)
  binary_mux_s1_w1 \picorv32_core/mux21_b9  (
    .i0(\picorv32_core/n57 [9]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n58 ),
    .o(\picorv32_core/n59 [9]));  // ../src/picorv32.v(449)
  binary_mux_s1_w1 \picorv32_core/mux22_b0  (
    .i0(\picorv32_core/n59 [0]),
    .i1(\picorv32_core/n68 [0]),
    .sel(\picorv32_core/n203 ),
    .o(\picorv32_core/n69 [0]));  // ../src/picorv32.v(456)
  binary_mux_s1_w1 \picorv32_core/mux22_b1  (
    .i0(\picorv32_core/n59 [1]),
    .i1(\picorv32_core/n68 [1]),
    .sel(\picorv32_core/n203 ),
    .o(\picorv32_core/n69 [1]));  // ../src/picorv32.v(456)
  binary_mux_s1_w1 \picorv32_core/mux22_b2  (
    .i0(\picorv32_core/n59 [2]),
    .i1(\picorv32_core/n68 [2]),
    .sel(\picorv32_core/n203 ),
    .o(\picorv32_core/n69 [2]));  // ../src/picorv32.v(456)
  binary_mux_s1_w1 \picorv32_core/mux22_b3  (
    .i0(\picorv32_core/n59 [3]),
    .i1(1'b0),
    .sel(\picorv32_core/n203 ),
    .o(\picorv32_core/n69 [3]));  // ../src/picorv32.v(456)
  binary_mux_s1_w1 \picorv32_core/mux22_b4  (
    .i0(\picorv32_core/n59 [4]),
    .i1(1'b0),
    .sel(\picorv32_core/n203 ),
    .o(\picorv32_core/n69 [4]));  // ../src/picorv32.v(456)
  binary_mux_s1_w1 \picorv32_core/mux22_b5  (
    .i0(\picorv32_core/n59 [5]),
    .i1(1'b0),
    .sel(\picorv32_core/n203 ),
    .o(\picorv32_core/n69 [5]));  // ../src/picorv32.v(456)
  binary_mux_s1_w1 \picorv32_core/mux22_b6  (
    .i0(\picorv32_core/n59 [6]),
    .i1(1'b0),
    .sel(\picorv32_core/n203 ),
    .o(\picorv32_core/n69 [6]));  // ../src/picorv32.v(456)
  binary_mux_s1_w1 \picorv32_core/mux22_b7  (
    .i0(\picorv32_core/n59 [7]),
    .i1(1'b0),
    .sel(\picorv32_core/n203 ),
    .o(\picorv32_core/n69 [7]));  // ../src/picorv32.v(456)
  binary_mux_s1_w1 \picorv32_core/mux22_b8  (
    .i0(\picorv32_core/n59 [8]),
    .i1(\picorv32_core/n61 ),
    .sel(\picorv32_core/n203 ),
    .o(\picorv32_core/n69 [8]));  // ../src/picorv32.v(456)
  binary_mux_s1_w1 \picorv32_core/mux22_b9  (
    .i0(\picorv32_core/n59 [9]),
    .i1(1'b0),
    .sel(\picorv32_core/n203 ),
    .o(\picorv32_core/n69 [9]));  // ../src/picorv32.v(456)
  binary_mux_s1_w1 \picorv32_core/mux23_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [2]),
    .sel(\picorv32_core/n99 ),
    .o(\picorv32_core/n192 [0]));  // ../src/picorv32.v(882)
  binary_mux_s1_w1 \picorv32_core/mux23_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [3]),
    .sel(\picorv32_core/n99 ),
    .o(\picorv32_core/n192 [1]));  // ../src/picorv32.v(882)
  binary_mux_s1_w1 \picorv32_core/mux23_b2  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [4]),
    .sel(\picorv32_core/n99 ),
    .o(\picorv32_core/n192 [2]));  // ../src/picorv32.v(882)
  binary_mux_s3_w1 \picorv32_core/mux24_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [12]),
    .i2(1'b0),
    .i3(\picorv32_core/n53 [0]),
    .i4(\picorv32_core/n69 [0]),
    .i5(\picorv32_core/n42 [12]),
    .i6(1'b0),
    .i7(1'b1),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [0]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [13]),
    .i2(1'b0),
    .i3(\picorv32_core/n53 [1]),
    .i4(\picorv32_core/n69 [1]),
    .i5(\picorv32_core/n42 [13]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [1]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b10  (
    .i0(\picorv32_core/mem_rdata_latched [4]),
    .i1(\picorv32_core/n42 [22]),
    .i2(\picorv32_core/mem_rdata_latched [4]),
    .i3(\picorv32_core/n53 [10]),
    .i4(\picorv32_core/n60 [2]),
    .i5(\picorv32_core/n42 [22]),
    .i6(\picorv32_core/n42 [22]),
    .i7(\picorv32_core/n42 [22]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [10]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b11  (
    .i0(\picorv32_core/mem_rdata_latched [5]),
    .i1(\picorv32_core/n42 [23]),
    .i2(\picorv32_core/mem_rdata_latched [5]),
    .i3(\picorv32_core/n53 [10]),
    .i4(\picorv32_core/n60 [3]),
    .i5(\picorv32_core/n42 [23]),
    .i6(\picorv32_core/n42 [23]),
    .i7(\picorv32_core/n42 [23]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [11]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b12  (
    .i0(\picorv32_core/mem_rdata_latched [6]),
    .i1(\picorv32_core/n42 [24]),
    .i2(\picorv32_core/mem_rdata_latched [6]),
    .i3(\picorv32_core/n53 [12]),
    .i4(\picorv32_core/n60 [4]),
    .i5(\picorv32_core/n42 [24]),
    .i6(\picorv32_core/n42 [24]),
    .i7(\picorv32_core/n42 [24]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [12]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b13  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/n42 [25]),
    .i2(\picorv32_core/mem_rdata_latched [12]),
    .i3(\picorv32_core/n53 [13]),
    .i4(\picorv32_core/n69 [3]),
    .i5(\picorv32_core/n42 [25]),
    .i6(\picorv32_core/mem_rdata_latched [2]),
    .i7(\picorv32_core/mem_rdata_latched [2]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [13]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b14  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/n42 [26]),
    .i2(\picorv32_core/mem_rdata_latched [12]),
    .i3(\picorv32_core/n53 [14]),
    .i4(\picorv32_core/n69 [4]),
    .i5(\picorv32_core/n42 [26]),
    .i6(\picorv32_core/mem_rdata_latched [5]),
    .i7(\picorv32_core/mem_rdata_latched [5]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [14]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b15  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/n42 [27]),
    .i2(\picorv32_core/mem_rdata_latched [12]),
    .i3(\picorv32_core/n53 [15]),
    .i4(\picorv32_core/n69 [5]),
    .i5(\picorv32_core/n42 [27]),
    .i6(\picorv32_core/mem_rdata_latched [6]),
    .i7(\picorv32_core/mem_rdata_latched [6]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [15]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b16  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/n42 [28]),
    .i2(\picorv32_core/mem_rdata_latched [12]),
    .i3(\picorv32_core/n53 [16]),
    .i4(\picorv32_core/n69 [6]),
    .i5(\picorv32_core/n42 [28]),
    .i6(\picorv32_core/mem_rdata_latched [12]),
    .i7(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [16]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b17  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/n42 [29]),
    .i2(\picorv32_core/mem_rdata_latched [12]),
    .i3(\picorv32_core/mem_rdata_latched [12]),
    .i4(\picorv32_core/n69 [7]),
    .i5(\picorv32_core/n42 [29]),
    .i6(\picorv32_core/mem_rdata_latched [12]),
    .i7(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [17]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b18  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/n42 [30]),
    .i2(\picorv32_core/mem_rdata_latched [12]),
    .i3(\picorv32_core/mem_rdata_latched [12]),
    .i4(\picorv32_core/n69 [8]),
    .i5(\picorv32_core/n42 [30]),
    .i6(\picorv32_core/mem_rdata_latched [12]),
    .i7(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [18]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b19  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/n42 [31]),
    .i2(\picorv32_core/mem_rdata_latched [12]),
    .i3(\picorv32_core/mem_rdata_latched [12]),
    .i4(\picorv32_core/n69 [9]),
    .i5(\picorv32_core/n42 [31]),
    .i6(\picorv32_core/mem_rdata_latched [12]),
    .i7(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [19]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b2  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [14]),
    .i2(1'b0),
    .i3(\picorv32_core/n53 [2]),
    .i4(\picorv32_core/n69 [2]),
    .i5(\picorv32_core/n42 [14]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [2]));  // ../src/picorv32.v(470)
  and \picorv32_core/mux24_b3_sel_is_3  (\picorv32_core/mux24_b3_sel_is_3_o , \picorv32_core/mem_rdata_latched [13], \picorv32_core/mem_rdata_latched [14], \picorv32_core/mem_rdata_latched$15$_neg , \picorv32_core/n193_neg );
  binary_mux_s3_w1 \picorv32_core/mux24_b8  (
    .i0(\picorv32_core/mem_rdata_latched [2]),
    .i1(\picorv32_core/n42 [20]),
    .i2(\picorv32_core/mem_rdata_latched [2]),
    .i3(\picorv32_core/n53 [10]),
    .i4(\picorv32_core/n60 [0]),
    .i5(\picorv32_core/n42 [20]),
    .i6(\picorv32_core/n42 [20]),
    .i7(\picorv32_core/n42 [20]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [8]));  // ../src/picorv32.v(470)
  binary_mux_s3_w1 \picorv32_core/mux24_b9  (
    .i0(\picorv32_core/mem_rdata_latched [3]),
    .i1(\picorv32_core/n42 [21]),
    .i2(\picorv32_core/mem_rdata_latched [3]),
    .i3(\picorv32_core/n53 [10]),
    .i4(\picorv32_core/n60 [1]),
    .i5(\picorv32_core/n42 [21]),
    .i6(\picorv32_core/n42 [21]),
    .i7(\picorv32_core/n42 [21]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n70 [9]));  // ../src/picorv32.v(470)
  and \picorv32_core/mux28_b0_sel_is_0  (\picorv32_core/mux28_b0_sel_is_0_o , \picorv32_core/n80_neg , \picorv32_core/n74_neg );
  binary_mux_s1_w1 \picorv32_core/mux2_b0  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [0]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [16]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [0]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b1  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [1]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [17]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [1]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b10  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [10]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [26]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [10]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b11  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [11]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [27]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [11]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b12  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [12]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [28]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [12]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b13  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [13]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [29]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [13]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b14  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [14]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [30]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [14]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b15  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [15]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [31]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [15]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b2  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [2]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [18]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [2]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b3  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [3]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [19]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [3]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b4  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [4]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [20]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [4]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b5  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [5]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [21]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [5]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b6  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [6]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [22]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [6]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b7  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [7]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [23]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [7]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b8  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [8]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [24]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [8]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux2_b9  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [9]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [25]),
    .sel(\picorv32_core/mem_la_firstword ),
    .o(\picorv32_core/n31 [9]));  // ../src/picorv32.v(352)
  and \picorv32_core/mux32_b0_sel_is_2  (\picorv32_core/mux32_b0_sel_is_2_o , \picorv32_core/n87_neg , \picorv32_core/mux28_b0_sel_is_0_o );
  AL_MUX \picorv32_core/mux35_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [14]),
    .sel(\picorv32_core/mux35_b0_sel_is_2_o ),
    .o(\picorv32_core/n93 [0]));
  and \picorv32_core/mux35_b0_sel_is_2  (\picorv32_core/mux35_b0_sel_is_2_o , \picorv32_core/n92_neg , \picorv32_core/mux32_b0_sel_is_2_o );
  AL_MUX \picorv32_core/mux35_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [28]),
    .sel(\picorv32_core/mux35_b0_sel_is_2_o ),
    .o(\picorv32_core/n93 [1]));
  AL_MUX \picorv32_core/mux35_b2  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [29]),
    .sel(\picorv32_core/mux35_b0_sel_is_2_o ),
    .o(\picorv32_core/n93 [2]));
  AL_MUX \picorv32_core/mux35_b3  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [30]),
    .sel(\picorv32_core/mux35_b0_sel_is_2_o ),
    .o(\picorv32_core/n93 [3]));
  AL_MUX \picorv32_core/mux35_b4  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [31]),
    .sel(\picorv32_core/mux35_b0_sel_is_2_o ),
    .o(\picorv32_core/n93 [4]));
  AL_MUX \picorv32_core/mux36_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [26]),
    .sel(\picorv32_core/mux35_b0_sel_is_2_o ),
    .o(\picorv32_core/n94 [0]));
  AL_MUX \picorv32_core/mux36_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [27]),
    .sel(\picorv32_core/mux35_b0_sel_is_2_o ),
    .o(\picorv32_core/n94 [1]));
  AL_MUX \picorv32_core/mux37_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [12]),
    .sel(\picorv32_core/mux35_b0_sel_is_2_o ),
    .o(\picorv32_core/n95 [0]));
  AL_MUX \picorv32_core/mux37_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [13]),
    .sel(\picorv32_core/mux35_b0_sel_is_2_o ),
    .o(\picorv32_core/n95 [1]));
  AL_MUX \picorv32_core/mux37_b2  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [25]),
    .sel(\picorv32_core/mux35_b0_sel_is_2_o ),
    .o(\picorv32_core/n95 [2]));
  AL_MUX \picorv32_core/mux38_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [20]),
    .sel(\picorv32_core/mux38_b0_sel_is_0_o ),
    .o(\picorv32_core/n91 [0]));
  and \picorv32_core/mux38_b0_sel_is_0  (\picorv32_core/mux38_b0_sel_is_0_o , \picorv32_core/n87_neg , \picorv32_core/n74_neg );
  AL_MUX \picorv32_core/mux38_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [21]),
    .sel(\picorv32_core/mux38_b0_sel_is_0_o ),
    .o(\picorv32_core/n91 [1]));
  AL_MUX \picorv32_core/mux38_b2  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [22]),
    .sel(\picorv32_core/mux38_b0_sel_is_0_o ),
    .o(\picorv32_core/n91 [2]));
  AL_MUX \picorv32_core/mux38_b3  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [23]),
    .sel(\picorv32_core/mux38_b0_sel_is_0_o ),
    .o(\picorv32_core/n91 [3]));
  AL_MUX \picorv32_core/mux38_b4  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [24]),
    .sel(\picorv32_core/mux38_b0_sel_is_0_o ),
    .o(\picorv32_core/n91 [4]));
  binary_mux_s1_w1 \picorv32_core/mux39_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [12]),
    .sel(\picorv32_core/n44 ),
    .o(\picorv32_core/n45 [0]));  // ../src/picorv32.v(416)
  binary_mux_s1_w1 \picorv32_core/mux39_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [14]),
    .sel(\picorv32_core/n44 ),
    .o(\picorv32_core/n45 [1]));  // ../src/picorv32.v(416)
  binary_mux_s1_w1 \picorv32_core/mux39_b2  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(\picorv32_core/n42 [25]),
    .sel(\picorv32_core/n44 ),
    .o(\picorv32_core/n45 [2]));  // ../src/picorv32.v(416)
  binary_mux_s1_w1 \picorv32_core/mux39_b3  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [30]),
    .sel(\picorv32_core/n44 ),
    .o(\picorv32_core/n45 [3]));  // ../src/picorv32.v(416)
  binary_mux_s1_w1 \picorv32_core/mux39_b4  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [31]),
    .sel(\picorv32_core/n44 ),
    .o(\picorv32_core/n45 [4]));  // ../src/picorv32.v(416)
  AL_MUX \picorv32_core/mux3_b16  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [0]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [16]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [16]));
  and \picorv32_core/mux3_b16_sel_is_0  (\picorv32_core/mux3_b16_sel_is_0_o , \picorv32_core/mem_la_secondword_neg , \picorv32_core/mem_la_firstword_neg );
  AL_MUX \picorv32_core/mux3_b17  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [1]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [17]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [17]));
  AL_MUX \picorv32_core/mux3_b18  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [2]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [18]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [18]));
  AL_MUX \picorv32_core/mux3_b19  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [3]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [19]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [19]));
  AL_MUX \picorv32_core/mux3_b20  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [4]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [20]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [20]));
  AL_MUX \picorv32_core/mux3_b21  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [5]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [21]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [21]));
  AL_MUX \picorv32_core/mux3_b22  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [6]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [22]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [22]));
  AL_MUX \picorv32_core/mux3_b23  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [7]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [23]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [23]));
  AL_MUX \picorv32_core/mux3_b24  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [8]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [24]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [24]));
  AL_MUX \picorv32_core/mux3_b25  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [9]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [25]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [25]));
  AL_MUX \picorv32_core/mux3_b26  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [10]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [26]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [26]));
  AL_MUX \picorv32_core/mux3_b27  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [11]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [27]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [27]));
  AL_MUX \picorv32_core/mux3_b28  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [12]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [28]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [28]));
  AL_MUX \picorv32_core/mux3_b29  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [13]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [29]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [29]));
  AL_MUX \picorv32_core/mux3_b30  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [14]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [30]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [30]));
  AL_MUX \picorv32_core/mux3_b31  (
    .i0(\picorv32_core/mem_rdata_latched_noshuffle [15]),
    .i1(\picorv32_core/mem_rdata_latched_noshuffle [31]),
    .sel(\picorv32_core/mux3_b16_sel_is_0_o ),
    .o(\picorv32_core/n32 [31]));
  binary_mux_s1_w1 \picorv32_core/mux40_b0  (
    .i0(\picorv32_core/n42 [20]),
    .i1(1'b0),
    .sel(\picorv32_core/n188 ),
    .o(\picorv32_core/n49 [0]));  // ../src/picorv32.v(416)
  binary_mux_s1_w1 \picorv32_core/mux40_b1  (
    .i0(\picorv32_core/n42 [21]),
    .i1(1'b0),
    .sel(\picorv32_core/n188 ),
    .o(\picorv32_core/n49 [1]));  // ../src/picorv32.v(416)
  binary_mux_s1_w1 \picorv32_core/mux40_b2  (
    .i0(\picorv32_core/n42 [22]),
    .i1(\picorv32_core/mem_rdata_latched [6]),
    .sel(\picorv32_core/n188 ),
    .o(\picorv32_core/n49 [2]));  // ../src/picorv32.v(416)
  binary_mux_s1_w1 \picorv32_core/mux40_b3  (
    .i0(\picorv32_core/n42 [24]),
    .i1(\picorv32_core/mem_rdata_latched [11]),
    .sel(\picorv32_core/n188 ),
    .o(\picorv32_core/n49 [3]));  // ../src/picorv32.v(416)
  binary_mux_s2_w1 \picorv32_core/mux41_b0  (
    .i0(\picorv32_core/n52 [0]),
    .i1(\picorv32_core/n71 [0]),
    .i2(\picorv32_core/n52 [0]),
    .i3(\picorv32_core/n42 [7]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [0]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b1  (
    .i0(\picorv32_core/n52 [1]),
    .i1(\picorv32_core/n71 [1]),
    .i2(\picorv32_core/n52 [1]),
    .i3(\picorv32_core/n42 [8]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [1]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b13  (
    .i0(\picorv32_core/n49 [0]),
    .i1(\picorv32_core/n70 [8]),
    .i2(\picorv32_core/n107 [0]),
    .i3(\picorv32_core/n42 [20]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [13]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b14  (
    .i0(\picorv32_core/n49 [1]),
    .i1(\picorv32_core/n70 [9]),
    .i2(\picorv32_core/n107 [1]),
    .i3(\picorv32_core/n42 [21]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [14]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b15  (
    .i0(\picorv32_core/n49 [2]),
    .i1(\picorv32_core/n70 [10]),
    .i2(\picorv32_core/n107 [2]),
    .i3(\picorv32_core/n42 [22]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [15]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b16  (
    .i0(\picorv32_core/n51 ),
    .i1(\picorv32_core/n70 [11]),
    .i2(\picorv32_core/n107 [3]),
    .i3(\picorv32_core/n42 [23]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [16]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b17  (
    .i0(\picorv32_core/n49 [3]),
    .i1(\picorv32_core/n70 [12]),
    .i2(\picorv32_core/n107 [4]),
    .i3(\picorv32_core/n42 [24]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [17]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b18  (
    .i0(\picorv32_core/n45 [2]),
    .i1(\picorv32_core/n70 [13]),
    .i2(\picorv32_core/n105 [2]),
    .i3(\picorv32_core/n42 [25]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [18]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b19  (
    .i0(\picorv32_core/n47 [1]),
    .i1(\picorv32_core/n70 [14]),
    .i2(\picorv32_core/n103 [0]),
    .i3(\picorv32_core/n42 [26]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [19]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b2  (
    .i0(\picorv32_core/n52 [2]),
    .i1(\picorv32_core/n71 [2]),
    .i2(\picorv32_core/n108 [2]),
    .i3(\picorv32_core/n42 [9]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [2]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b20  (
    .i0(\picorv32_core/n47 [2]),
    .i1(\picorv32_core/n70 [15]),
    .i2(\picorv32_core/n103 [1]),
    .i3(\picorv32_core/n42 [27]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [20]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b21  (
    .i0(\picorv32_core/n47 [3]),
    .i1(\picorv32_core/n70 [16]),
    .i2(\picorv32_core/n102 [1]),
    .i3(\picorv32_core/n42 [28]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [21]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b22  (
    .i0(\picorv32_core/n47 [4]),
    .i1(\picorv32_core/n70 [17]),
    .i2(\picorv32_core/n102 [2]),
    .i3(\picorv32_core/n42 [29]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [22]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b23  (
    .i0(\picorv32_core/n45 [3]),
    .i1(\picorv32_core/n70 [18]),
    .i2(\picorv32_core/n102 [3]),
    .i3(\picorv32_core/n42 [30]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [23]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b24  (
    .i0(\picorv32_core/n45 [4]),
    .i1(\picorv32_core/n70 [19]),
    .i2(\picorv32_core/n102 [4]),
    .i3(\picorv32_core/n42 [31]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [24]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b3  (
    .i0(\picorv32_core/n52 [3]),
    .i1(\picorv32_core/n71 [3]),
    .i2(\picorv32_core/n52 [3]),
    .i3(\picorv32_core/n42 [10]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [3]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b4  (
    .i0(\picorv32_core/n52 [4]),
    .i1(\picorv32_core/n71 [4]),
    .i2(\picorv32_core/n52 [4]),
    .i3(\picorv32_core/n42 [11]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [4]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b5  (
    .i0(\picorv32_core/n45 [0]),
    .i1(\picorv32_core/n70 [0]),
    .i2(\picorv32_core/n105 [0]),
    .i3(\picorv32_core/n42 [12]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [5]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b6  (
    .i0(\picorv32_core/n47 [0]),
    .i1(\picorv32_core/n70 [1]),
    .i2(\picorv32_core/n105 [1]),
    .i3(\picorv32_core/n42 [13]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [6]));  // ../src/picorv32.v(506)
  binary_mux_s2_w1 \picorv32_core/mux41_b7  (
    .i0(\picorv32_core/n45 [1]),
    .i1(\picorv32_core/n70 [2]),
    .i2(\picorv32_core/n102 [0]),
    .i3(\picorv32_core/n42 [14]),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n109 [7]));  // ../src/picorv32.v(506)
  binary_mux_s1_w1 \picorv32_core/mux42_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_state [0]),
    .sel(resetn),
    .o(\picorv32_core/n112 [0]));  // ../src/picorv32.v(532)
  binary_mux_s1_w1 \picorv32_core/mux42_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_state [1]),
    .sel(resetn),
    .o(\picorv32_core/n112 [1]));  // ../src/picorv32.v(532)
  binary_mux_s1_w1 \picorv32_core/mux47_b0  (
    .i0(\picorv32_core/mem_state [0]),
    .i1(1'b1),
    .sel(\picorv32_core/n120 ),
    .o(\picorv32_core/n124 [0]));  // ../src/picorv32.v(552)
  binary_mux_s1_w1 \picorv32_core/mux47_b1  (
    .i0(\picorv32_core/mem_state [1]),
    .i1(1'b0),
    .sel(\picorv32_core/n120 ),
    .o(\picorv32_core/n124 [1]));  // ../src/picorv32.v(552)
  binary_mux_s1_w1 \picorv32_core/mux48_b0  (
    .i0(\picorv32_core/n124 [0]),
    .i1(1'b0),
    .sel(\picorv32_core/mem_do_wdata ),
    .o(\picorv32_core/n127 [0]));  // ../src/picorv32.v(557)
  binary_mux_s1_w1 \picorv32_core/mux48_b1  (
    .i0(\picorv32_core/n124 [1]),
    .i1(1'b1),
    .sel(\picorv32_core/mem_do_wdata ),
    .o(\picorv32_core/n127 [1]));  // ../src/picorv32.v(557)
  binary_mux_s1_w1 \picorv32_core/mux49_b0  (
    .i0(mem_rdata[16]),
    .i1(\picorv32_core/mem_16bit_buffer [0]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [0]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b1  (
    .i0(mem_rdata[17]),
    .i1(\picorv32_core/mem_16bit_buffer [1]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [1]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b10  (
    .i0(mem_rdata[26]),
    .i1(\picorv32_core/mem_16bit_buffer [10]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [10]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b11  (
    .i0(mem_rdata[27]),
    .i1(\picorv32_core/mem_16bit_buffer [11]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [11]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b12  (
    .i0(mem_rdata[28]),
    .i1(\picorv32_core/mem_16bit_buffer [12]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [12]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b13  (
    .i0(mem_rdata[29]),
    .i1(\picorv32_core/mem_16bit_buffer [13]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [13]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b14  (
    .i0(mem_rdata[30]),
    .i1(\picorv32_core/mem_16bit_buffer [14]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [14]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b15  (
    .i0(mem_rdata[31]),
    .i1(\picorv32_core/mem_16bit_buffer [15]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [15]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b2  (
    .i0(mem_rdata[18]),
    .i1(\picorv32_core/mem_16bit_buffer [2]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [2]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b3  (
    .i0(mem_rdata[19]),
    .i1(\picorv32_core/mem_16bit_buffer [3]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [3]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b4  (
    .i0(mem_rdata[20]),
    .i1(\picorv32_core/mem_16bit_buffer [4]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [4]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b5  (
    .i0(mem_rdata[21]),
    .i1(\picorv32_core/mem_16bit_buffer [5]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [5]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b6  (
    .i0(mem_rdata[22]),
    .i1(\picorv32_core/mem_16bit_buffer [6]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [6]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b7  (
    .i0(mem_rdata[23]),
    .i1(\picorv32_core/mem_16bit_buffer [7]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [7]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b8  (
    .i0(mem_rdata[24]),
    .i1(\picorv32_core/mem_16bit_buffer [8]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [8]));  // ../src/picorv32.v(569)
  binary_mux_s1_w1 \picorv32_core/mux49_b9  (
    .i0(mem_rdata[25]),
    .i1(\picorv32_core/mem_16bit_buffer [9]),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/n128 [9]));  // ../src/picorv32.v(569)
  AL_MUX \picorv32_core/mux4_b0  (
    .i0(\picorv32_core/mem_16bit_buffer [0]),
    .i1(\picorv32_core/n31 [0]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [0]));
  and \picorv32_core/mux4_b0_sel_is_0  (\picorv32_core/mux4_b0_sel_is_0_o , \picorv32_core/mem_la_use_prefetched_high_word_neg , \picorv32_core/mem_la_secondword_neg );
  AL_MUX \picorv32_core/mux4_b1  (
    .i0(\picorv32_core/mem_16bit_buffer [1]),
    .i1(\picorv32_core/n31 [1]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [1]));
  AL_MUX \picorv32_core/mux4_b10  (
    .i0(\picorv32_core/mem_16bit_buffer [10]),
    .i1(\picorv32_core/n31 [10]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [10]));
  AL_MUX \picorv32_core/mux4_b11  (
    .i0(\picorv32_core/mem_16bit_buffer [11]),
    .i1(\picorv32_core/n31 [11]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [11]));
  AL_MUX \picorv32_core/mux4_b12  (
    .i0(\picorv32_core/mem_16bit_buffer [12]),
    .i1(\picorv32_core/n31 [12]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [12]));
  AL_MUX \picorv32_core/mux4_b13  (
    .i0(\picorv32_core/mem_16bit_buffer [13]),
    .i1(\picorv32_core/n31 [13]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [13]));
  AL_MUX \picorv32_core/mux4_b14  (
    .i0(\picorv32_core/mem_16bit_buffer [14]),
    .i1(\picorv32_core/n31 [14]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [14]));
  AL_MUX \picorv32_core/mux4_b15  (
    .i0(\picorv32_core/mem_16bit_buffer [15]),
    .i1(\picorv32_core/n31 [15]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [15]));
  binary_mux_s1_w1 \picorv32_core/mux4_b16  (
    .i0(\picorv32_core/n32 [16]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [16]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b17  (
    .i0(\picorv32_core/n32 [17]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [17]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b18  (
    .i0(\picorv32_core/n32 [18]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [18]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b19  (
    .i0(\picorv32_core/n32 [19]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [19]));  // ../src/picorv32.v(352)
  AL_MUX \picorv32_core/mux4_b2  (
    .i0(\picorv32_core/mem_16bit_buffer [2]),
    .i1(\picorv32_core/n31 [2]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [2]));
  binary_mux_s1_w1 \picorv32_core/mux4_b20  (
    .i0(\picorv32_core/n32 [20]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [20]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b21  (
    .i0(\picorv32_core/n32 [21]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [21]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b22  (
    .i0(\picorv32_core/n32 [22]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [22]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b23  (
    .i0(\picorv32_core/n32 [23]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [23]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b24  (
    .i0(\picorv32_core/n32 [24]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [24]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b25  (
    .i0(\picorv32_core/n32 [25]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [25]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b26  (
    .i0(\picorv32_core/n32 [26]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [26]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b27  (
    .i0(\picorv32_core/n32 [27]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [27]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b28  (
    .i0(\picorv32_core/n32 [28]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [28]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b29  (
    .i0(\picorv32_core/n32 [29]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [29]));  // ../src/picorv32.v(352)
  AL_MUX \picorv32_core/mux4_b3  (
    .i0(\picorv32_core/mem_16bit_buffer [3]),
    .i1(\picorv32_core/n31 [3]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [3]));
  binary_mux_s1_w1 \picorv32_core/mux4_b30  (
    .i0(\picorv32_core/n32 [30]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [30]));  // ../src/picorv32.v(352)
  binary_mux_s1_w1 \picorv32_core/mux4_b31  (
    .i0(\picorv32_core/n32 [31]),
    .i1(1'bx),
    .sel(\picorv32_core/mem_la_use_prefetched_high_word ),
    .o(\picorv32_core/mem_rdata_latched [31]));  // ../src/picorv32.v(352)
  AL_MUX \picorv32_core/mux4_b4  (
    .i0(\picorv32_core/mem_16bit_buffer [4]),
    .i1(\picorv32_core/n31 [4]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [4]));
  AL_MUX \picorv32_core/mux4_b5  (
    .i0(\picorv32_core/mem_16bit_buffer [5]),
    .i1(\picorv32_core/n31 [5]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [5]));
  AL_MUX \picorv32_core/mux4_b6  (
    .i0(\picorv32_core/mem_16bit_buffer [6]),
    .i1(\picorv32_core/n31 [6]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [6]));
  AL_MUX \picorv32_core/mux4_b7  (
    .i0(\picorv32_core/mem_16bit_buffer [7]),
    .i1(\picorv32_core/n31 [7]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [7]));
  AL_MUX \picorv32_core/mux4_b8  (
    .i0(\picorv32_core/mem_16bit_buffer [8]),
    .i1(\picorv32_core/n31 [8]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [8]));
  AL_MUX \picorv32_core/mux4_b9  (
    .i0(\picorv32_core/mem_16bit_buffer [9]),
    .i1(\picorv32_core/n31 [9]),
    .sel(\picorv32_core/mux4_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_latched [9]));
  AL_MUX \picorv32_core/mux51_b0  (
    .i0(\picorv32_core/mem_16bit_buffer [0]),
    .i1(mem_rdata[16]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [0]));
  and \picorv32_core/mux51_b0_sel_is_3  (\picorv32_core/mux51_b0_sel_is_3_o , \picorv32_core/n598 , \picorv32_core/n131 );
  AL_MUX \picorv32_core/mux51_b1  (
    .i0(\picorv32_core/mem_16bit_buffer [1]),
    .i1(mem_rdata[17]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [1]));
  AL_MUX \picorv32_core/mux51_b10  (
    .i0(\picorv32_core/mem_16bit_buffer [10]),
    .i1(mem_rdata[26]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [10]));
  AL_MUX \picorv32_core/mux51_b11  (
    .i0(\picorv32_core/mem_16bit_buffer [11]),
    .i1(mem_rdata[27]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [11]));
  AL_MUX \picorv32_core/mux51_b12  (
    .i0(\picorv32_core/mem_16bit_buffer [12]),
    .i1(mem_rdata[28]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [12]));
  AL_MUX \picorv32_core/mux51_b13  (
    .i0(\picorv32_core/mem_16bit_buffer [13]),
    .i1(mem_rdata[29]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [13]));
  AL_MUX \picorv32_core/mux51_b14  (
    .i0(\picorv32_core/mem_16bit_buffer [14]),
    .i1(mem_rdata[30]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [14]));
  AL_MUX \picorv32_core/mux51_b15  (
    .i0(\picorv32_core/mem_16bit_buffer [15]),
    .i1(mem_rdata[31]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [15]));
  AL_MUX \picorv32_core/mux51_b2  (
    .i0(\picorv32_core/mem_16bit_buffer [2]),
    .i1(mem_rdata[18]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [2]));
  AL_MUX \picorv32_core/mux51_b3  (
    .i0(\picorv32_core/mem_16bit_buffer [3]),
    .i1(mem_rdata[19]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [3]));
  AL_MUX \picorv32_core/mux51_b4  (
    .i0(\picorv32_core/mem_16bit_buffer [4]),
    .i1(mem_rdata[20]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [4]));
  AL_MUX \picorv32_core/mux51_b5  (
    .i0(\picorv32_core/mem_16bit_buffer [5]),
    .i1(mem_rdata[21]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [5]));
  AL_MUX \picorv32_core/mux51_b6  (
    .i0(\picorv32_core/mem_16bit_buffer [6]),
    .i1(mem_rdata[22]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [6]));
  AL_MUX \picorv32_core/mux51_b7  (
    .i0(\picorv32_core/mem_16bit_buffer [7]),
    .i1(mem_rdata[23]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [7]));
  AL_MUX \picorv32_core/mux51_b8  (
    .i0(\picorv32_core/mem_16bit_buffer [8]),
    .i1(mem_rdata[24]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [8]));
  AL_MUX \picorv32_core/mux51_b9  (
    .i0(\picorv32_core/mem_16bit_buffer [9]),
    .i1(mem_rdata[25]),
    .sel(\picorv32_core/mux51_b0_sel_is_3_o ),
    .o(\picorv32_core/n133 [9]));
  binary_mux_s1_w1 \picorv32_core/mux52_b0  (
    .i0(\picorv32_core/n133 [0]),
    .i1(\picorv32_core/n128 [0]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [0]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b1  (
    .i0(\picorv32_core/n133 [1]),
    .i1(\picorv32_core/n128 [1]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [1]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b10  (
    .i0(\picorv32_core/n133 [10]),
    .i1(\picorv32_core/n128 [10]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [10]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b11  (
    .i0(\picorv32_core/n133 [11]),
    .i1(\picorv32_core/n128 [11]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [11]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b12  (
    .i0(\picorv32_core/n133 [12]),
    .i1(\picorv32_core/n128 [12]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [12]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b13  (
    .i0(\picorv32_core/n133 [13]),
    .i1(\picorv32_core/n128 [13]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [13]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b14  (
    .i0(\picorv32_core/n133 [14]),
    .i1(\picorv32_core/n128 [14]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [14]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b15  (
    .i0(\picorv32_core/n133 [15]),
    .i1(\picorv32_core/n128 [15]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [15]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b2  (
    .i0(\picorv32_core/n133 [2]),
    .i1(\picorv32_core/n128 [2]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [2]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b3  (
    .i0(\picorv32_core/n133 [3]),
    .i1(\picorv32_core/n128 [3]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [3]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b4  (
    .i0(\picorv32_core/n133 [4]),
    .i1(\picorv32_core/n128 [4]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [4]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b5  (
    .i0(\picorv32_core/n133 [5]),
    .i1(\picorv32_core/n128 [5]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [5]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b6  (
    .i0(\picorv32_core/n133 [6]),
    .i1(\picorv32_core/n128 [6]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [6]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b7  (
    .i0(\picorv32_core/n133 [7]),
    .i1(\picorv32_core/n128 [7]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [7]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b8  (
    .i0(\picorv32_core/n133 [8]),
    .i1(\picorv32_core/n128 [8]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [8]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux52_b9  (
    .i0(\picorv32_core/n133 [9]),
    .i1(\picorv32_core/n128 [9]),
    .sel(\picorv32_core/mem_la_read ),
    .o(\picorv32_core/n136 [9]));  // ../src/picorv32.v(582)
  binary_mux_s1_w1 \picorv32_core/mux55_b0  (
    .i0(\picorv32_core/n42 [7]),
    .i1(\picorv32_core/n109 [0]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [0]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b1  (
    .i0(\picorv32_core/n42 [8]),
    .i1(\picorv32_core/n109 [1]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [1]));  // ../src/picorv32.v(507)
  AL_MUX \picorv32_core/mux55_b10  (
    .i0(\picorv32_core/n42 [17]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/mux55_b10_sel_is_3_o ),
    .o(\picorv32_core/n110 [10]));
  and \picorv32_core/mux55_b10_sel_is_3  (\picorv32_core/mux55_b10_sel_is_3_o , \picorv32_core/n43 , \picorv32_core/mux105_sel_is_5_o );
  AL_MUX \picorv32_core/mux55_b11  (
    .i0(\picorv32_core/n42 [18]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/mux55_b10_sel_is_3_o ),
    .o(\picorv32_core/n110 [11]));
  AL_MUX \picorv32_core/mux55_b12  (
    .i0(\picorv32_core/n42 [19]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/mux55_b10_sel_is_3_o ),
    .o(\picorv32_core/n110 [12]));
  binary_mux_s1_w1 \picorv32_core/mux55_b13  (
    .i0(\picorv32_core/n42 [20]),
    .i1(\picorv32_core/n109 [13]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [13]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b14  (
    .i0(\picorv32_core/n42 [21]),
    .i1(\picorv32_core/n109 [14]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [14]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b15  (
    .i0(\picorv32_core/n42 [22]),
    .i1(\picorv32_core/n109 [15]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [15]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b16  (
    .i0(\picorv32_core/n42 [23]),
    .i1(\picorv32_core/n109 [16]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [16]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b17  (
    .i0(\picorv32_core/n42 [24]),
    .i1(\picorv32_core/n109 [17]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [17]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b18  (
    .i0(\picorv32_core/n42 [25]),
    .i1(\picorv32_core/n109 [18]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [18]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b19  (
    .i0(\picorv32_core/n42 [26]),
    .i1(\picorv32_core/n109 [19]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [19]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b2  (
    .i0(\picorv32_core/n42 [9]),
    .i1(\picorv32_core/n109 [2]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [2]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b20  (
    .i0(\picorv32_core/n42 [27]),
    .i1(\picorv32_core/n109 [20]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [20]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b21  (
    .i0(\picorv32_core/n42 [28]),
    .i1(\picorv32_core/n109 [21]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [21]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b22  (
    .i0(\picorv32_core/n42 [29]),
    .i1(\picorv32_core/n109 [22]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [22]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b23  (
    .i0(\picorv32_core/n42 [30]),
    .i1(\picorv32_core/n109 [23]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [23]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b24  (
    .i0(\picorv32_core/n42 [31]),
    .i1(\picorv32_core/n109 [24]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [24]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b3  (
    .i0(\picorv32_core/n42 [10]),
    .i1(\picorv32_core/n109 [3]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [3]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b4  (
    .i0(\picorv32_core/n42 [11]),
    .i1(\picorv32_core/n109 [4]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [4]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b5  (
    .i0(\picorv32_core/n42 [12]),
    .i1(\picorv32_core/n109 [5]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [5]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b6  (
    .i0(\picorv32_core/n42 [13]),
    .i1(\picorv32_core/n109 [6]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [6]));  // ../src/picorv32.v(507)
  binary_mux_s1_w1 \picorv32_core/mux55_b7  (
    .i0(\picorv32_core/n42 [14]),
    .i1(\picorv32_core/n109 [7]),
    .sel(\picorv32_core/n43 ),
    .o(\picorv32_core/n110 [7]));  // ../src/picorv32.v(507)
  AL_MUX \picorv32_core/mux55_b8  (
    .i0(\picorv32_core/n42 [15]),
    .i1(\picorv32_core/mem_rdata_latched [5]),
    .sel(\picorv32_core/mux55_b10_sel_is_3_o ),
    .o(\picorv32_core/n110 [8]));
  AL_MUX \picorv32_core/mux55_b9  (
    .i0(\picorv32_core/n42 [16]),
    .i1(\picorv32_core/mem_rdata_latched [6]),
    .sel(\picorv32_core/mux55_b10_sel_is_3_o ),
    .o(\picorv32_core/n110 [9]));
  binary_mux_s1_w1 \picorv32_core/mux56_b0  (
    .i0(\picorv32_core/mem_state [0]),
    .i1(1'b0),
    .sel(\picorv32_core/mem_do_rinst ),
    .o(\picorv32_core/n146 [0]));  // ../src/picorv32.v(598)
  binary_mux_s1_w1 \picorv32_core/mux56_b1  (
    .i0(\picorv32_core/mem_state [1]),
    .i1(1'b0),
    .sel(\picorv32_core/mem_do_rinst ),
    .o(\picorv32_core/n146 [1]));  // ../src/picorv32.v(598)
  binary_mux_s2_w1 \picorv32_core/mux57_b0  (
    .i0(\picorv32_core/n127 [0]),
    .i1(\picorv32_core/n143 [0]),
    .i2(\picorv32_core/n145 [0]),
    .i3(\picorv32_core/n146 [0]),
    .sel(\picorv32_core/mem_state ),
    .o(\picorv32_core/n147 [0]));  // ../src/picorv32.v(600)
  binary_mux_s2_w1 \picorv32_core/mux57_b1  (
    .i0(\picorv32_core/n127 [1]),
    .i1(\picorv32_core/n143 [1]),
    .i2(\picorv32_core/n145 [1]),
    .i3(\picorv32_core/n146 [1]),
    .sel(\picorv32_core/mem_state ),
    .o(\picorv32_core/n147 [1]));  // ../src/picorv32.v(600)
  binary_mux_s2_w1 \picorv32_core/mux58  (
    .i0(\picorv32_core/n125 ),
    .i1(\picorv32_core/n139 ),
    .i2(\picorv32_core/n144 ),
    .i3(\picorv32_core/mem_valid ),
    .sel(\picorv32_core/mem_state ),
    .o(\picorv32_core/n148 ));  // ../src/picorv32.v(600)
  and \picorv32_core/mux59_sel_is_5  (\picorv32_core/mux59_sel_is_5_o , \picorv32_core/mem_state [0], \picorv32_core/mem_state$1$_neg , \picorv32_core/mem_xfer );
  binary_mux_s1_w1 \picorv32_core/mux5_b0  (
    .i0(mem_rdata[0]),
    .i1(mem_rdata[16]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [0]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b1  (
    .i0(mem_rdata[1]),
    .i1(mem_rdata[17]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [1]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b10  (
    .i0(mem_rdata[10]),
    .i1(mem_rdata[26]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [10]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b11  (
    .i0(mem_rdata[11]),
    .i1(mem_rdata[27]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [11]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b12  (
    .i0(mem_rdata[12]),
    .i1(mem_rdata[28]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [12]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b13  (
    .i0(mem_rdata[13]),
    .i1(mem_rdata[29]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [13]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b14  (
    .i0(mem_rdata[14]),
    .i1(mem_rdata[30]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [14]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b15  (
    .i0(mem_rdata[15]),
    .i1(mem_rdata[31]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [15]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b2  (
    .i0(mem_rdata[2]),
    .i1(mem_rdata[18]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [2]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b3  (
    .i0(mem_rdata[3]),
    .i1(mem_rdata[19]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [3]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b4  (
    .i0(mem_rdata[4]),
    .i1(mem_rdata[20]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [4]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b5  (
    .i0(mem_rdata[5]),
    .i1(mem_rdata[21]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [5]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b6  (
    .i0(mem_rdata[6]),
    .i1(mem_rdata[22]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [6]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b7  (
    .i0(mem_rdata[7]),
    .i1(mem_rdata[23]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [7]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b8  (
    .i0(mem_rdata[8]),
    .i1(mem_rdata[24]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [8]));  // ../src/picorv32.v(379)
  binary_mux_s1_w1 \picorv32_core/mux5_b9  (
    .i0(mem_rdata[9]),
    .i1(mem_rdata[25]),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n39 [9]));  // ../src/picorv32.v(379)
  and \picorv32_core/mux61_sel_is_5  (\picorv32_core/mux61_sel_is_5_o , \picorv32_core/mem_state [0], \picorv32_core/mem_state$1$_neg , \picorv32_core/u173_sel_is_3_o );
  binary_mux_s1_w1 \picorv32_core/mux64_b0  (
    .i0(\picorv32_core/n147 [0]),
    .i1(\picorv32_core/n112 [0]),
    .sel(\picorv32_core/n111 ),
    .o(\picorv32_core/n154 [0]));  // ../src/picorv32.v(601)
  binary_mux_s1_w1 \picorv32_core/mux64_b1  (
    .i0(\picorv32_core/n147 [1]),
    .i1(\picorv32_core/n112 [1]),
    .sel(\picorv32_core/n111 ),
    .o(\picorv32_core/n154 [1]));  // ../src/picorv32.v(601)
  and \picorv32_core/mux68_b0_sel_is_2  (\picorv32_core/mux68_b0_sel_is_2_o , \picorv32_core/n111_neg , \picorv32_core/mux59_sel_is_5_o );
  AL_MUX \picorv32_core/mux69_b0  (
    .i0(\picorv32_core/mem_state [0]),
    .i1(\picorv32_core/n135 [0]),
    .sel(\picorv32_core/mux69_b0_sel_is_1_o ),
    .o(\picorv32_core/n143 [0]));
  and \picorv32_core/mux69_b0_sel_is_1  (\picorv32_core/mux69_b0_sel_is_1_o , \picorv32_core/mem_xfer , \picorv32_core/mem_la_read_neg );
  AL_MUX \picorv32_core/mux69_b1  (
    .i0(\picorv32_core/mem_state [1]),
    .i1(\picorv32_core/n135 [0]),
    .sel(\picorv32_core/mux69_b0_sel_is_1_o ),
    .o(\picorv32_core/n143 [1]));
  binary_mux_s1_w1 \picorv32_core/mux69_b2  (
    .i0(\picorv32_core/mem_state [0]),
    .i1(1'b0),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n145 [0]));  // ../src/picorv32.v(591)
  binary_mux_s1_w1 \picorv32_core/mux69_b3  (
    .i0(\picorv32_core/mem_state [1]),
    .i1(1'b0),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n145 [1]));  // ../src/picorv32.v(591)
  binary_mux_s2_w1 \picorv32_core/mux6_b0  (
    .i0(mem_rdata[0]),
    .i1(mem_rdata[8]),
    .i2(mem_rdata[16]),
    .i3(mem_rdata[24]),
    .sel({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .o(\picorv32_core/n41 [0]));  // ../src/picorv32.v(389)
  binary_mux_s2_w1 \picorv32_core/mux6_b1  (
    .i0(mem_rdata[1]),
    .i1(mem_rdata[9]),
    .i2(mem_rdata[17]),
    .i3(mem_rdata[25]),
    .sel({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .o(\picorv32_core/n41 [1]));  // ../src/picorv32.v(389)
  binary_mux_s2_w1 \picorv32_core/mux6_b2  (
    .i0(mem_rdata[2]),
    .i1(mem_rdata[10]),
    .i2(mem_rdata[18]),
    .i3(mem_rdata[26]),
    .sel({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .o(\picorv32_core/n41 [2]));  // ../src/picorv32.v(389)
  binary_mux_s2_w1 \picorv32_core/mux6_b3  (
    .i0(mem_rdata[3]),
    .i1(mem_rdata[11]),
    .i2(mem_rdata[19]),
    .i3(mem_rdata[27]),
    .sel({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .o(\picorv32_core/n41 [3]));  // ../src/picorv32.v(389)
  binary_mux_s2_w1 \picorv32_core/mux6_b4  (
    .i0(mem_rdata[4]),
    .i1(mem_rdata[12]),
    .i2(mem_rdata[20]),
    .i3(mem_rdata[28]),
    .sel({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .o(\picorv32_core/n41 [4]));  // ../src/picorv32.v(389)
  binary_mux_s2_w1 \picorv32_core/mux6_b5  (
    .i0(mem_rdata[5]),
    .i1(mem_rdata[13]),
    .i2(mem_rdata[21]),
    .i3(mem_rdata[29]),
    .sel({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .o(\picorv32_core/n41 [5]));  // ../src/picorv32.v(389)
  binary_mux_s2_w1 \picorv32_core/mux6_b6  (
    .i0(mem_rdata[6]),
    .i1(mem_rdata[14]),
    .i2(mem_rdata[22]),
    .i3(mem_rdata[30]),
    .sel({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .o(\picorv32_core/n41 [6]));  // ../src/picorv32.v(389)
  binary_mux_s2_w1 \picorv32_core/mux6_b7  (
    .i0(mem_rdata[7]),
    .i1(mem_rdata[15]),
    .i2(mem_rdata[23]),
    .i3(mem_rdata[31]),
    .sel({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .o(\picorv32_core/n41 [7]));  // ../src/picorv32.v(389)
  binary_mux_s1_w1 \picorv32_core/mux70_b0  (
    .i0(\picorv32_core/mem_rdata_latched [7]),
    .i1(1'b0),
    .sel(\picorv32_core/n184 ),
    .o(\picorv32_core/n186 [0]));  // ../src/picorv32.v(882)
  binary_mux_s1_w1 \picorv32_core/mux70_b1  (
    .i0(\picorv32_core/mem_rdata_latched [9]),
    .i1(1'b0),
    .sel(\picorv32_core/n184 ),
    .o(\picorv32_core/n186 [1]));  // ../src/picorv32.v(882)
  binary_mux_s1_w1 \picorv32_core/mux71_b0  (
    .i0(\picorv32_core/mem_rdata_latched [21]),
    .i1(\picorv32_core/mem_rdata_latched [3]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [0]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b1  (
    .i0(\picorv32_core/mem_rdata_latched [22]),
    .i1(\picorv32_core/mem_rdata_latched [4]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [1]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b10  (
    .i0(\picorv32_core/mem_rdata_latched [20]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [10]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b11  (
    .i0(\picorv32_core/mem_rdata_latched [13]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [11]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b12  (
    .i0(\picorv32_core/mem_rdata_latched [14]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [12]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b13  (
    .i0(\picorv32_core/mem_rdata_latched [15]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [13]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b14  (
    .i0(\picorv32_core/mem_rdata_latched [16]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [14]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b15  (
    .i0(\picorv32_core/mem_rdata_latched [17]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [15]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b16  (
    .i0(\picorv32_core/mem_rdata_latched [18]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [16]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b17  (
    .i0(\picorv32_core/mem_rdata_latched [19]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [17]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b18  (
    .i0(\picorv32_core/mem_rdata_latched [31]),
    .i1(\picorv32_core/mem_rdata_latched [12]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [18]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b2  (
    .i0(\picorv32_core/mem_rdata_latched [23]),
    .i1(\picorv32_core/mem_rdata_latched [5]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [2]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b3  (
    .i0(\picorv32_core/mem_rdata_latched [24]),
    .i1(\picorv32_core/mem_rdata_latched [11]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [3]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b4  (
    .i0(\picorv32_core/mem_rdata_latched [25]),
    .i1(\picorv32_core/mem_rdata_latched [2]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [4]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b5  (
    .i0(\picorv32_core/mem_rdata_latched [26]),
    .i1(\picorv32_core/mem_rdata_latched [7]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [5]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b6  (
    .i0(\picorv32_core/mem_rdata_latched [27]),
    .i1(\picorv32_core/mem_rdata_latched [6]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [6]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b7  (
    .i0(\picorv32_core/mem_rdata_latched [28]),
    .i1(\picorv32_core/mem_rdata_latched [9]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [7]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b8  (
    .i0(\picorv32_core/mem_rdata_latched [29]),
    .i1(\picorv32_core/mem_rdata_latched [10]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [8]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux71_b9  (
    .i0(\picorv32_core/mem_rdata_latched [30]),
    .i1(\picorv32_core/mem_rdata_latched [8]),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n248 [9]));  // ../src/picorv32.v(990)
  binary_mux_s1_w1 \picorv32_core/mux72_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [7]),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n195 [0]));  // ../src/picorv32.v(909)
  binary_mux_s1_w1 \picorv32_core/mux72_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [8]),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n195 [1]));  // ../src/picorv32.v(909)
  binary_mux_s1_w1 \picorv32_core/mux72_b2  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [9]),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n195 [2]));  // ../src/picorv32.v(909)
  binary_mux_s1_w1 \picorv32_core/mux72_b3  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [10]),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n195 [3]));  // ../src/picorv32.v(909)
  binary_mux_s1_w1 \picorv32_core/mux72_b4  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [11]),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n195 [4]));  // ../src/picorv32.v(909)
  binary_mux_s1_w1 \picorv32_core/mux74_b3  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [5]),
    .sel(\picorv32_core/n197 ),
    .o(\picorv32_core/n200 [3]));  // ../src/picorv32.v(917)
  and \picorv32_core/mux75_b0_sel_is_0  (\picorv32_core/mux75_b0_sel_is_0_o , \picorv32_core/n58_neg , \picorv32_core/mem_rdata_latched [11]);
  AL_MUX \picorv32_core/mux76_b0  (
    .i0(\picorv32_core/mem_rdata_latched [7]),
    .i1(1'b0),
    .sel(\picorv32_core/mux76_b0_sel_is_2_o ),
    .o(\picorv32_core/n205 [0]));
  and \picorv32_core/mux76_b0_sel_is_2  (\picorv32_core/mux76_b0_sel_is_2_o , \picorv32_core/n203_neg , \picorv32_core/mux75_b0_sel_is_0_o );
  AL_MUX \picorv32_core/mux76_b1  (
    .i0(\picorv32_core/mem_rdata_latched [8]),
    .i1(1'b0),
    .sel(\picorv32_core/mux76_b0_sel_is_2_o ),
    .o(\picorv32_core/n205 [1]));
  AL_MUX \picorv32_core/mux76_b2  (
    .i0(\picorv32_core/mem_rdata_latched [9]),
    .i1(1'b0),
    .sel(\picorv32_core/mux76_b0_sel_is_2_o ),
    .o(\picorv32_core/n205 [2]));
  AL_MUX \picorv32_core/mux76_b3  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\picorv32_core/mux76_b0_sel_is_2_o ),
    .o(\picorv32_core/n205 [3]));
  and \picorv32_core/mux77_b0_sel_is_0  (\picorv32_core/mux77_b0_sel_is_0_o , \picorv32_core/n203_neg , \picorv32_core/mem_rdata_latched [11]);
  not \picorv32_core/mux77_b0_sel_is_0_o_inv  (\picorv32_core/mux77_b0_sel_is_0_o_neg , \picorv32_core/mux77_b0_sel_is_0_o );
  binary_mux_s1_w1 \picorv32_core/mux77_b3  (
    .i0(\picorv32_core/n200 [3]),
    .i1(1'b1),
    .sel(\picorv32_core/n203 ),
    .o(\picorv32_core/n206 [3]));  // ../src/picorv32.v(928)
  and \picorv32_core/mux77_b4_sel_is_2  (\picorv32_core/mux77_b4_sel_is_2_o , \picorv32_core/n203_neg , \picorv32_core/n197 );
  binary_mux_s3_w1 \picorv32_core/mux79_b0  (
    .i0(\picorv32_core/mem_rdata_latched [7]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(\picorv32_core/n195 [0]),
    .i4(\picorv32_core/n205 [0]),
    .i5(1'b0),
    .i6(\picorv32_core/mem_rdata_latched [7]),
    .i7(\picorv32_core/mem_rdata_latched [7]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n208 [0]));  // ../src/picorv32.v(943)
  binary_mux_s3_w1 \picorv32_core/mux79_b1  (
    .i0(\picorv32_core/mem_rdata_latched [8]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(\picorv32_core/n195 [1]),
    .i4(\picorv32_core/n205 [1]),
    .i5(1'b0),
    .i6(\picorv32_core/mem_rdata_latched [8]),
    .i7(\picorv32_core/mem_rdata_latched [8]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n208 [1]));  // ../src/picorv32.v(943)
  binary_mux_s3_w1 \picorv32_core/mux79_b2  (
    .i0(\picorv32_core/mem_rdata_latched [9]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(\picorv32_core/n195 [2]),
    .i4(\picorv32_core/n205 [2]),
    .i5(1'b0),
    .i6(\picorv32_core/mem_rdata_latched [9]),
    .i7(\picorv32_core/mem_rdata_latched [9]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n208 [2]));  // ../src/picorv32.v(943)
  binary_mux_s3_w1 \picorv32_core/mux79_b3  (
    .i0(\picorv32_core/mem_rdata_latched [10]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(\picorv32_core/n195 [3]),
    .i4(\picorv32_core/n205 [3]),
    .i5(1'b0),
    .i6(1'b1),
    .i7(1'b1),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n208 [3]));  // ../src/picorv32.v(943)
  binary_mux_s3_w1 \picorv32_core/mux79_b4  (
    .i0(\picorv32_core/mem_rdata_latched [11]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(\picorv32_core/n195 [4]),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n208 [4]));  // ../src/picorv32.v(943)
  binary_mux_s1_w1 \picorv32_core/mux7_b0  (
    .i0(\picorv32_core/pcpi_rs2$8$ ),
    .i1(mem_la_wdata[0]),
    .sel(\picorv32_core/mem_wordsize [1]),
    .o(mem_la_wdata[8]));  // ../src/picorv32.v(391)
  binary_mux_s1_w1 \picorv32_core/mux7_b1  (
    .i0(\picorv32_core/pcpi_rs2$9$ ),
    .i1(mem_la_wdata[1]),
    .sel(\picorv32_core/mem_wordsize [1]),
    .o(mem_la_wdata[9]));  // ../src/picorv32.v(391)
  binary_mux_s1_w1 \picorv32_core/mux7_b2  (
    .i0(\picorv32_core/pcpi_rs2$10$ ),
    .i1(mem_la_wdata[2]),
    .sel(\picorv32_core/mem_wordsize [1]),
    .o(mem_la_wdata[10]));  // ../src/picorv32.v(391)
  binary_mux_s1_w1 \picorv32_core/mux7_b3  (
    .i0(\picorv32_core/pcpi_rs2$11$ ),
    .i1(mem_la_wdata[3]),
    .sel(\picorv32_core/mem_wordsize [1]),
    .o(mem_la_wdata[11]));  // ../src/picorv32.v(391)
  binary_mux_s1_w1 \picorv32_core/mux7_b4  (
    .i0(\picorv32_core/pcpi_rs2$12$ ),
    .i1(mem_la_wdata[4]),
    .sel(\picorv32_core/mem_wordsize [1]),
    .o(mem_la_wdata[12]));  // ../src/picorv32.v(391)
  binary_mux_s1_w1 \picorv32_core/mux7_b5  (
    .i0(\picorv32_core/pcpi_rs2$13$ ),
    .i1(mem_la_wdata[5]),
    .sel(\picorv32_core/mem_wordsize [1]),
    .o(mem_la_wdata[13]));  // ../src/picorv32.v(391)
  binary_mux_s1_w1 \picorv32_core/mux7_b6  (
    .i0(\picorv32_core/pcpi_rs2$14$ ),
    .i1(mem_la_wdata[6]),
    .sel(\picorv32_core/mem_wordsize [1]),
    .o(mem_la_wdata[14]));  // ../src/picorv32.v(391)
  binary_mux_s1_w1 \picorv32_core/mux7_b7  (
    .i0(\picorv32_core/pcpi_rs2$15$ ),
    .i1(mem_la_wdata[7]),
    .sel(\picorv32_core/mem_wordsize [1]),
    .o(mem_la_wdata[15]));  // ../src/picorv32.v(391)
  AL_MUX \picorv32_core/mux80_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [2]),
    .sel(\picorv32_core/mux80_b0_sel_is_4_o ),
    .o(\picorv32_core/n209 [0]));
  and \picorv32_core/mux80_b0_sel_is_4  (\picorv32_core/mux80_b0_sel_is_4_o , \picorv32_core/mem_rdata_latched$13$_neg , \picorv32_core/mem_rdata_latched$14$_neg , \picorv32_core/mem_rdata_latched [15], \picorv32_core/mux77_b0_sel_is_0_o_neg );
  AL_MUX \picorv32_core/mux80_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [3]),
    .sel(\picorv32_core/mux80_b0_sel_is_4_o ),
    .o(\picorv32_core/n209 [1]));
  AL_MUX \picorv32_core/mux80_b2  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [4]),
    .sel(\picorv32_core/mux80_b0_sel_is_4_o ),
    .o(\picorv32_core/n209 [2]));
  AL_MUX \picorv32_core/mux80_b3  (
    .i0(1'b0),
    .i1(\picorv32_core/n206 [3]),
    .sel(\picorv32_core/mux80_b3_sel_is_4_o ),
    .o(\picorv32_core/n209 [3]));
  and \picorv32_core/mux80_b3_sel_is_4  (\picorv32_core/mux80_b3_sel_is_4_o , \picorv32_core/mem_rdata_latched$13$_neg , \picorv32_core/mem_rdata_latched$14$_neg , \picorv32_core/mem_rdata_latched [15]);
  AL_MUX \picorv32_core/mux80_b4  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [6]),
    .sel(\picorv32_core/mux80_b4_sel_is_12_o ),
    .o(\picorv32_core/n209 [4]));
  and \picorv32_core/mux80_b4_sel_is_12  (\picorv32_core/mux80_b4_sel_is_12_o , \picorv32_core/mem_rdata_latched$13$_neg , \picorv32_core/mem_rdata_latched$14$_neg , \picorv32_core/mem_rdata_latched [15], \picorv32_core/mux77_b4_sel_is_2_o );
  and \picorv32_core/mux81_sel_is_1  (\picorv32_core/mux81_sel_is_1_o , \picorv32_core/mem_rdata_latched [13], \picorv32_core/mem_rdata_latched$14$_neg );
  binary_mux_s3_w1 \picorv32_core/mux82  (
    .i0(1'b1),
    .i1(\picorv32_core/n178 ),
    .i2(1'b1),
    .i3(\picorv32_core/n194 ),
    .i4(\picorv32_core/n201 ),
    .i5(\picorv32_core/n178 ),
    .i6(\picorv32_core/n178 ),
    .i7(\picorv32_core/n178 ),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n211 ));  // ../src/picorv32.v(943)
  binary_mux_s3_w1 \picorv32_core/mux83_b0  (
    .i0(\picorv32_core/mem_rdata_latched [7]),
    .i1(1'b1),
    .i2(\picorv32_core/mem_rdata_latched [7]),
    .i3(\picorv32_core/mem_rdata_latched [7]),
    .i4(\picorv32_core/n205 [0]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n212 [0]));  // ../src/picorv32.v(943)
  binary_mux_s3_w1 \picorv32_core/mux83_b1  (
    .i0(\picorv32_core/mem_rdata_latched [8]),
    .i1(1'b0),
    .i2(\picorv32_core/mem_rdata_latched [8]),
    .i3(\picorv32_core/mem_rdata_latched [8]),
    .i4(\picorv32_core/n205 [1]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n212 [1]));  // ../src/picorv32.v(943)
  binary_mux_s3_w1 \picorv32_core/mux83_b2  (
    .i0(\picorv32_core/mem_rdata_latched [9]),
    .i1(1'b0),
    .i2(\picorv32_core/mem_rdata_latched [9]),
    .i3(\picorv32_core/mem_rdata_latched [9]),
    .i4(\picorv32_core/n205 [2]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n212 [2]));  // ../src/picorv32.v(943)
  binary_mux_s3_w1 \picorv32_core/mux83_b3  (
    .i0(\picorv32_core/mem_rdata_latched [10]),
    .i1(1'b0),
    .i2(\picorv32_core/mem_rdata_latched [10]),
    .i3(\picorv32_core/mem_rdata_latched [10]),
    .i4(\picorv32_core/n205 [3]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n212 [3]));  // ../src/picorv32.v(943)
  binary_mux_s3_w1 \picorv32_core/mux83_b4  (
    .i0(\picorv32_core/mem_rdata_latched [11]),
    .i1(1'b0),
    .i2(\picorv32_core/mem_rdata_latched [11]),
    .i3(\picorv32_core/mem_rdata_latched [11]),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n212 [4]));  // ../src/picorv32.v(943)
  AL_MUX \picorv32_core/mux84  (
    .i0(\picorv32_core/n179 ),
    .i1(1'b1),
    .sel(\picorv32_core/mux84_sel_is_12_o ),
    .o(\picorv32_core/n213 ));
  and \picorv32_core/mux84_sel_is_12  (\picorv32_core/mux84_sel_is_12_o , \picorv32_core/mem_rdata_latched$13$_neg , \picorv32_core/mem_rdata_latched$14$_neg , \picorv32_core/mem_rdata_latched [15], \picorv32_core/n203 );
  binary_mux_s1_w1 \picorv32_core/mux87_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/mem_rdata_latched [7]),
    .sel(\picorv32_core/n80 ),
    .o(\picorv32_core/n218 [0]));  // ../src/picorv32.v(969)
  and \picorv32_core/mux88_b0_sel_is_2  (\picorv32_core/mux88_b0_sel_is_2_o , \picorv32_core/n80_neg , \picorv32_core/n74 );
  not \picorv32_core/mux88_b0_sel_is_2_o_inv  (\picorv32_core/mux88_b0_sel_is_2_o_neg , \picorv32_core/mux88_b0_sel_is_2_o );
  binary_mux_s2_w1 \picorv32_core/mux8_b0  (
    .i0(1'b1),
    .i1(\picorv32_core/n38 [0]),
    .i2(\picorv32_core/n40 [0]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(mem_la_wstrb[0]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux8_b1  (
    .i0(1'b1),
    .i1(\picorv32_core/n38 [0]),
    .i2(\picorv32_core/n40 [1]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(mem_la_wstrb[1]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux8_b2  (
    .i0(1'b1),
    .i1(\picorv32_core/pcpi_rs1$1$ ),
    .i2(\picorv32_core/n40 [2]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(mem_la_wstrb[2]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux8_b3  (
    .i0(1'b1),
    .i1(\picorv32_core/pcpi_rs1$1$ ),
    .i2(\picorv32_core/n40 [3]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(mem_la_wstrb[3]));  // ../src/picorv32.v(391)
  binary_mux_s1_w1 \picorv32_core/mux90_b0  (
    .i0(\picorv32_core/n218 [0]),
    .i1(1'b1),
    .sel(\picorv32_core/n87 ),
    .o(\picorv32_core/n222 [0]));  // ../src/picorv32.v(974)
  and \picorv32_core/mux90_b1_sel_is_2  (\picorv32_core/mux90_b1_sel_is_2_o , \picorv32_core/n87_neg , \picorv32_core/n80 );
  not \picorv32_core/mux90_b1_sel_is_2_o_inv  (\picorv32_core/mux90_b1_sel_is_2_o_neg , \picorv32_core/mux90_b1_sel_is_2_o );
  and \picorv32_core/mux91_b0_sel_is_0  (\picorv32_core/mux91_b0_sel_is_0_o , \picorv32_core/n87_neg , \picorv32_core/mux88_b0_sel_is_2_o_neg );
  binary_mux_s1_w1 \picorv32_core/mux92_b0  (
    .i0(\picorv32_core/n222 [0]),
    .i1(\picorv32_core/mem_rdata_latched [7]),
    .sel(\picorv32_core/n92 ),
    .o(\picorv32_core/n225 [0]));  // ../src/picorv32.v(980)
  AL_MUX \picorv32_core/mux92_b1  (
    .i0(\picorv32_core/mem_rdata_latched [8]),
    .i1(1'b0),
    .sel(\picorv32_core/mux92_b1_sel_is_0_o ),
    .o(\picorv32_core/n225 [1]));
  and \picorv32_core/mux92_b1_sel_is_0  (\picorv32_core/mux92_b1_sel_is_0_o , \picorv32_core/n92_neg , \picorv32_core/mux90_b1_sel_is_2_o_neg );
  AL_MUX \picorv32_core/mux92_b2  (
    .i0(\picorv32_core/mem_rdata_latched [9]),
    .i1(1'b0),
    .sel(\picorv32_core/mux92_b1_sel_is_0_o ),
    .o(\picorv32_core/n225 [2]));
  AL_MUX \picorv32_core/mux92_b3  (
    .i0(\picorv32_core/mem_rdata_latched [10]),
    .i1(1'b0),
    .sel(\picorv32_core/mux92_b1_sel_is_0_o ),
    .o(\picorv32_core/n225 [3]));
  AL_MUX \picorv32_core/mux92_b4  (
    .i0(\picorv32_core/mem_rdata_latched [11]),
    .i1(1'b0),
    .sel(\picorv32_core/mux92_b1_sel_is_0_o ),
    .o(\picorv32_core/n225 [4]));
  AL_MUX \picorv32_core/mux93_b0  (
    .i0(\picorv32_core/mem_rdata_latched [7]),
    .i1(1'b0),
    .sel(\picorv32_core/mux93_b0_sel_is_2_o ),
    .o(\picorv32_core/n226 [0]));
  and \picorv32_core/mux93_b0_sel_is_2  (\picorv32_core/mux93_b0_sel_is_2_o , \picorv32_core/n92_neg , \picorv32_core/mux91_b0_sel_is_0_o );
  AL_MUX \picorv32_core/mux93_b1  (
    .i0(\picorv32_core/mem_rdata_latched [8]),
    .i1(1'b0),
    .sel(\picorv32_core/mux93_b0_sel_is_2_o ),
    .o(\picorv32_core/n226 [1]));
  AL_MUX \picorv32_core/mux93_b2  (
    .i0(\picorv32_core/mem_rdata_latched [9]),
    .i1(1'b0),
    .sel(\picorv32_core/mux93_b0_sel_is_2_o ),
    .o(\picorv32_core/n226 [2]));
  AL_MUX \picorv32_core/mux93_b3  (
    .i0(\picorv32_core/mem_rdata_latched [10]),
    .i1(1'b0),
    .sel(\picorv32_core/mux93_b0_sel_is_2_o ),
    .o(\picorv32_core/n226 [3]));
  AL_MUX \picorv32_core/mux93_b4  (
    .i0(\picorv32_core/mem_rdata_latched [11]),
    .i1(1'b0),
    .sel(\picorv32_core/mux93_b0_sel_is_2_o ),
    .o(\picorv32_core/n226 [4]));
  AL_MUX \picorv32_core/mux94_b0  (
    .i0(\picorv32_core/mem_rdata_latched [2]),
    .i1(1'b0),
    .sel(\picorv32_core/mux94_b0_sel_is_0_o ),
    .o(\picorv32_core/n227 [0]));
  and \picorv32_core/mux94_b0_sel_is_0  (\picorv32_core/mux94_b0_sel_is_0_o , \picorv32_core/n92_neg , \picorv32_core/n80_neg );
  AL_MUX \picorv32_core/mux94_b1  (
    .i0(\picorv32_core/mem_rdata_latched [3]),
    .i1(1'b0),
    .sel(\picorv32_core/mux94_b0_sel_is_0_o ),
    .o(\picorv32_core/n227 [1]));
  AL_MUX \picorv32_core/mux94_b2  (
    .i0(\picorv32_core/mem_rdata_latched [4]),
    .i1(1'b0),
    .sel(\picorv32_core/mux94_b0_sel_is_0_o ),
    .o(\picorv32_core/n227 [2]));
  AL_MUX \picorv32_core/mux94_b3  (
    .i0(\picorv32_core/mem_rdata_latched [5]),
    .i1(1'b0),
    .sel(\picorv32_core/mux94_b0_sel_is_0_o ),
    .o(\picorv32_core/n227 [3]));
  AL_MUX \picorv32_core/mux94_b4  (
    .i0(\picorv32_core/mem_rdata_latched [6]),
    .i1(1'b0),
    .sel(\picorv32_core/mux94_b0_sel_is_0_o ),
    .o(\picorv32_core/n227 [4]));
  binary_mux_s2_w1 \picorv32_core/mux95  (
    .i0(\picorv32_core/n183 ),
    .i1(\picorv32_core/n211 ),
    .i2(\picorv32_core/n228 ),
    .i3(\picorv32_core/n178 ),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n234 ));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux96_b0  (
    .i0(\picorv32_core/n189 [0]),
    .i1(\picorv32_core/n212 [0]),
    .i2(\picorv32_core/n229 [0]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n235 [0]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux96_b1  (
    .i0(\picorv32_core/n189 [1]),
    .i1(\picorv32_core/n212 [1]),
    .i2(\picorv32_core/n229 [1]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n235 [1]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux96_b2  (
    .i0(\picorv32_core/n189 [2]),
    .i1(\picorv32_core/n212 [2]),
    .i2(\picorv32_core/n229 [2]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n235 [2]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux96_b3  (
    .i0(\picorv32_core/n188 ),
    .i1(\picorv32_core/n212 [3]),
    .i2(\picorv32_core/n229 [3]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n235 [3]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux96_b4  (
    .i0(1'b0),
    .i1(\picorv32_core/n212 [4]),
    .i2(\picorv32_core/n229 [4]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n235 [4]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux97_b0  (
    .i0(\picorv32_core/n186 [0]),
    .i1(\picorv32_core/n208 [0]),
    .i2(\picorv32_core/n230 [0]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n236 [0]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux97_b1  (
    .i0(\picorv32_core/sel7/or_B1_B2_o ),
    .i1(\picorv32_core/n208 [1]),
    .i2(\picorv32_core/n230 [1]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n236 [1]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux97_b2  (
    .i0(\picorv32_core/n186 [1]),
    .i1(\picorv32_core/n208 [2]),
    .i2(\picorv32_core/n230 [2]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n236 [2]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux97_b3  (
    .i0(\picorv32_core/n185 ),
    .i1(\picorv32_core/n208 [3]),
    .i2(\picorv32_core/n230 [3]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n236 [3]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux97_b4  (
    .i0(1'b0),
    .i1(\picorv32_core/n208 [4]),
    .i2(\picorv32_core/n230 [4]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n236 [4]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux98_b0  (
    .i0(\picorv32_core/n192 [0]),
    .i1(\picorv32_core/n209 [0]),
    .i2(\picorv32_core/n231 [0]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n237 [0]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux98_b1  (
    .i0(\picorv32_core/n192 [1]),
    .i1(\picorv32_core/n209 [1]),
    .i2(\picorv32_core/n231 [1]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n237 [1]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux98_b2  (
    .i0(\picorv32_core/n192 [2]),
    .i1(\picorv32_core/n209 [2]),
    .i2(\picorv32_core/n231 [2]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n237 [2]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux98_b3  (
    .i0(\picorv32_core/n99 ),
    .i1(\picorv32_core/n209 [3]),
    .i2(\picorv32_core/n231 [3]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n237 [3]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux98_b4  (
    .i0(1'b0),
    .i1(\picorv32_core/n209 [4]),
    .i2(\picorv32_core/n231 [4]),
    .i3(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n237 [4]));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux99  (
    .i0(\picorv32_core/n190 ),
    .i1(\picorv32_core/n176 ),
    .i2(\picorv32_core/n190 ),
    .i3(\picorv32_core/n176 ),
    .sel(\picorv32_core/mem_rdata_latched [1:0]),
    .o(\picorv32_core/n238 ));  // ../src/picorv32.v(989)
  binary_mux_s2_w1 \picorv32_core/mux9_b0  (
    .i0(mem_rdata[0]),
    .i1(\picorv32_core/n39 [0]),
    .i2(\picorv32_core/n41 [0]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/n641 [0]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux9_b1  (
    .i0(mem_rdata[1]),
    .i1(\picorv32_core/n39 [1]),
    .i2(\picorv32_core/n41 [1]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/n641 [1]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux9_b10  (
    .i0(mem_rdata[10]),
    .i1(\picorv32_core/n39 [10]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/mem_rdata_word [10]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux9_b11  (
    .i0(mem_rdata[11]),
    .i1(\picorv32_core/n39 [11]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/mem_rdata_word [11]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux9_b12  (
    .i0(mem_rdata[12]),
    .i1(\picorv32_core/n39 [12]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/mem_rdata_word [12]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux9_b13  (
    .i0(mem_rdata[13]),
    .i1(\picorv32_core/n39 [13]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/mem_rdata_word [13]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux9_b14  (
    .i0(mem_rdata[14]),
    .i1(\picorv32_core/n39 [14]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/mem_rdata_word [14]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux9_b15  (
    .i0(mem_rdata[15]),
    .i1(\picorv32_core/n39 [15]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/mem_rdata_word [15]));  // ../src/picorv32.v(391)
  AL_MUX \picorv32_core/mux9_b16  (
    .i0(1'b0),
    .i1(mem_rdata[16]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [16]));
  AL_MUX \picorv32_core/mux9_b17  (
    .i0(1'b0),
    .i1(mem_rdata[17]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [17]));
  AL_MUX \picorv32_core/mux9_b18  (
    .i0(1'b0),
    .i1(mem_rdata[18]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [18]));
  AL_MUX \picorv32_core/mux9_b19  (
    .i0(1'b0),
    .i1(mem_rdata[19]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [19]));
  binary_mux_s2_w1 \picorv32_core/mux9_b2  (
    .i0(mem_rdata[2]),
    .i1(\picorv32_core/n39 [2]),
    .i2(\picorv32_core/n41 [2]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/n641 [2]));  // ../src/picorv32.v(391)
  AL_MUX \picorv32_core/mux9_b20  (
    .i0(1'b0),
    .i1(mem_rdata[20]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [20]));
  AL_MUX \picorv32_core/mux9_b21  (
    .i0(1'b0),
    .i1(mem_rdata[21]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [21]));
  AL_MUX \picorv32_core/mux9_b22  (
    .i0(1'b0),
    .i1(mem_rdata[22]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [22]));
  AL_MUX \picorv32_core/mux9_b23  (
    .i0(1'b0),
    .i1(mem_rdata[23]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [23]));
  AL_MUX \picorv32_core/mux9_b24  (
    .i0(1'b0),
    .i1(mem_rdata[24]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [24]));
  AL_MUX \picorv32_core/mux9_b25  (
    .i0(1'b0),
    .i1(mem_rdata[25]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [25]));
  AL_MUX \picorv32_core/mux9_b26  (
    .i0(1'b0),
    .i1(mem_rdata[26]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [26]));
  AL_MUX \picorv32_core/mux9_b27  (
    .i0(1'b0),
    .i1(mem_rdata[27]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [27]));
  AL_MUX \picorv32_core/mux9_b28  (
    .i0(1'b0),
    .i1(mem_rdata[28]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [28]));
  AL_MUX \picorv32_core/mux9_b29  (
    .i0(1'b0),
    .i1(mem_rdata[29]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [29]));
  binary_mux_s2_w1 \picorv32_core/mux9_b3  (
    .i0(mem_rdata[3]),
    .i1(\picorv32_core/n39 [3]),
    .i2(\picorv32_core/n41 [3]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/n641 [3]));  // ../src/picorv32.v(391)
  AL_MUX \picorv32_core/mux9_b30  (
    .i0(1'b0),
    .i1(mem_rdata[30]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [30]));
  AL_MUX \picorv32_core/mux9_b31  (
    .i0(1'b0),
    .i1(mem_rdata[31]),
    .sel(\picorv32_core/mux165_b0_sel_is_0_o ),
    .o(\picorv32_core/mem_rdata_word [31]));
  binary_mux_s2_w1 \picorv32_core/mux9_b4  (
    .i0(mem_rdata[4]),
    .i1(\picorv32_core/n39 [4]),
    .i2(\picorv32_core/n41 [4]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/n641 [4]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux9_b5  (
    .i0(mem_rdata[5]),
    .i1(\picorv32_core/n39 [5]),
    .i2(\picorv32_core/n41 [5]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/n641 [5]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux9_b6  (
    .i0(mem_rdata[6]),
    .i1(\picorv32_core/n39 [6]),
    .i2(\picorv32_core/n41 [6]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/n641 [6]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux9_b7  (
    .i0(mem_rdata[7]),
    .i1(\picorv32_core/n39 [7]),
    .i2(\picorv32_core/n41 [7]),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/n641 [7]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux9_b8  (
    .i0(mem_rdata[8]),
    .i1(\picorv32_core/n39 [8]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/mem_rdata_word [8]));  // ../src/picorv32.v(391)
  binary_mux_s2_w1 \picorv32_core/mux9_b9  (
    .i0(mem_rdata[9]),
    .i1(\picorv32_core/n39 [9]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\picorv32_core/mem_wordsize ),
    .o(\picorv32_core/mem_rdata_word [9]));  // ../src/picorv32.v(391)
  not \picorv32_core/n111_inv  (\picorv32_core/n111_neg , \picorv32_core/n111 );
  not \picorv32_core/n193_inv  (\picorv32_core/n193_neg , \picorv32_core/n193 );
  not \picorv32_core/n203_inv  (\picorv32_core/n203_neg , \picorv32_core/n203 );
  not \picorv32_core/n274_inv  (\picorv32_core/n274_neg , \picorv32_core/n274 );
  not \picorv32_core/n54_inv  (\picorv32_core/n54_neg , \picorv32_core/n54 );
  not \picorv32_core/n56_inv  (\picorv32_core/n56_neg , \picorv32_core/n56 );
  not \picorv32_core/n58_inv  (\picorv32_core/n58_neg , \picorv32_core/n58 );
  not \picorv32_core/n61_inv  (\picorv32_core/n61_neg , \picorv32_core/n61 );
  not \picorv32_core/n63_inv  (\picorv32_core/n63_neg , \picorv32_core/n63 );
  not \picorv32_core/n65_inv  (\picorv32_core/n65_neg , \picorv32_core/n65 );
  not \picorv32_core/n67_inv  (\picorv32_core/n67_neg , \picorv32_core/n67 );
  not \picorv32_core/n701_inv  (\picorv32_core/n701_neg , \picorv32_core/n701 );
  not \picorv32_core/n736_inv  (\picorv32_core/n736_neg , \picorv32_core/n736 );
  not \picorv32_core/n740_inv  (\picorv32_core/n740_neg , \picorv32_core/n740 );
  not \picorv32_core/n744_inv  (\picorv32_core/n744_neg , \picorv32_core/n744 );
  not \picorv32_core/n74_inv  (\picorv32_core/n74_neg , \picorv32_core/n74 );
  not \picorv32_core/n80_inv  (\picorv32_core/n80_neg , \picorv32_core/n80 );
  not \picorv32_core/n87_inv  (\picorv32_core/n87_neg , \picorv32_core/n87 );
  not \picorv32_core/n92_inv  (\picorv32_core/n92_neg , \picorv32_core/n92 );
  ne_w5 \picorv32_core/neq0  (
    .i0(\picorv32_core/mem_rdata_latched [6:2]),
    .i1(5'b00000),
    .o(\picorv32_core/n79 ));  // ../src/picorv32.v(487)
  ne_w1 \picorv32_core/neq1  (
    .i0(\picorv32_core/mem_rdata_latched [12]),
    .i1(1'b0),
    .o(\picorv32_core/n84 ));  // ../src/picorv32.v(491)
  ne_w5 \picorv32_core/neq2  (
    .i0(\picorv32_core/mem_rdata_latched [11:7]),
    .i1(5'b00000),
    .o(\picorv32_core/n85 ));  // ../src/picorv32.v(491)
  ne_w2 \picorv32_core/neq3  (
    .i0(\picorv32_core/mem_rdata_latched [1:0]),
    .i1(2'b11),
    .o(\picorv32_core/n180 ));  // ../src/picorv32.v(855)
  ne_w2 \picorv32_core/neq4  (
    .i0({\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .i1(2'b00),
    .o(\picorv32_core/n735 ));  // ../src/picorv32.v(1854)
  ne_w1 \picorv32_core/neq5  (
    .i0(\picorv32_core/pcpi_rs1$0$ ),
    .i1(1'b0),
    .o(\picorv32_core/n739 ));  // ../src/picorv32.v(1861)
  reg_sr_as_w1 \picorv32_core/prefetched_high_word_reg  (
    .clk(clk),
    .d(\picorv32_core/n131 ),
    .en(\picorv32_core/mux61_sel_is_5_o ),
    .reset(~\picorv32_core/u179_sel_is_0_o ),
    .set(1'b0),
    .q(\picorv32_core/prefetched_high_word ));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg0_b0  (
    .clk(clk),
    .d(\picorv32_core/mem_rdata_latched [0]),
    .en(\picorv32_core/mem_xfer ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [0]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b1  (
    .clk(clk),
    .d(\picorv32_core/mem_rdata_latched [1]),
    .en(\picorv32_core/mem_xfer ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [1]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b10  (
    .clk(clk),
    .d(\picorv32_core/n110 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [10]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b11  (
    .clk(clk),
    .d(\picorv32_core/n110 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [11]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b12  (
    .clk(clk),
    .d(\picorv32_core/n110 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [12]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b13  (
    .clk(clk),
    .d(\picorv32_core/n110 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [13]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b14  (
    .clk(clk),
    .d(\picorv32_core/n110 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [14]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b15  (
    .clk(clk),
    .d(\picorv32_core/n110 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [15]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b16  (
    .clk(clk),
    .d(\picorv32_core/n110 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [16]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b17  (
    .clk(clk),
    .d(\picorv32_core/n110 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [17]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b18  (
    .clk(clk),
    .d(\picorv32_core/n110 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [18]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b19  (
    .clk(clk),
    .d(\picorv32_core/n110 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [19]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b2  (
    .clk(clk),
    .d(\picorv32_core/mem_rdata_latched [2]),
    .en(\picorv32_core/mem_xfer ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [2]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b20  (
    .clk(clk),
    .d(\picorv32_core/n110 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [20]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b21  (
    .clk(clk),
    .d(\picorv32_core/n110 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [21]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b22  (
    .clk(clk),
    .d(\picorv32_core/n110 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [22]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b23  (
    .clk(clk),
    .d(\picorv32_core/n110 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [23]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b24  (
    .clk(clk),
    .d(\picorv32_core/n110 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [24]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b25  (
    .clk(clk),
    .d(\picorv32_core/n110 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [25]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b26  (
    .clk(clk),
    .d(\picorv32_core/n110 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [26]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b27  (
    .clk(clk),
    .d(\picorv32_core/n110 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [27]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b28  (
    .clk(clk),
    .d(\picorv32_core/n110 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [28]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b29  (
    .clk(clk),
    .d(\picorv32_core/n110 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [29]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b3  (
    .clk(clk),
    .d(\picorv32_core/mem_rdata_latched [3]),
    .en(\picorv32_core/mem_xfer ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [3]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b30  (
    .clk(clk),
    .d(\picorv32_core/n110 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [30]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b31  (
    .clk(clk),
    .d(\picorv32_core/n110 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [31]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b4  (
    .clk(clk),
    .d(\picorv32_core/mem_rdata_latched [4]),
    .en(\picorv32_core/mem_xfer ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [4]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b5  (
    .clk(clk),
    .d(\picorv32_core/mem_rdata_latched [5]),
    .en(\picorv32_core/mem_xfer ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [5]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b6  (
    .clk(clk),
    .d(\picorv32_core/mem_rdata_latched [6]),
    .en(\picorv32_core/mem_xfer ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [6]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b7  (
    .clk(clk),
    .d(\picorv32_core/n110 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [7]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b8  (
    .clk(clk),
    .d(\picorv32_core/n110 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [8]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg0_b9  (
    .clk(clk),
    .d(\picorv32_core/n110 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_rdata_q [9]));  // ../src/picorv32.v(508)
  reg_ar_as_w1 \picorv32_core/reg11_b0  (
    .clk(clk),
    .d(\picorv32_core/n358 [0]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [0]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b1  (
    .clk(clk),
    .d(\picorv32_core/n358 [1]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [1]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b10  (
    .clk(clk),
    .d(\picorv32_core/n358 [10]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [10]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b11  (
    .clk(clk),
    .d(\picorv32_core/n358 [11]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [11]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b12  (
    .clk(clk),
    .d(\picorv32_core/n358 [12]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [12]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b13  (
    .clk(clk),
    .d(\picorv32_core/n358 [13]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [13]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b14  (
    .clk(clk),
    .d(\picorv32_core/n358 [14]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [14]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b15  (
    .clk(clk),
    .d(\picorv32_core/n358 [15]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [15]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b16  (
    .clk(clk),
    .d(\picorv32_core/n358 [16]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [16]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b17  (
    .clk(clk),
    .d(\picorv32_core/n358 [17]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [17]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b18  (
    .clk(clk),
    .d(\picorv32_core/n358 [18]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [18]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b19  (
    .clk(clk),
    .d(\picorv32_core/n358 [19]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [19]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b2  (
    .clk(clk),
    .d(\picorv32_core/n358 [2]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [2]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b20  (
    .clk(clk),
    .d(\picorv32_core/n358 [20]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [20]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b21  (
    .clk(clk),
    .d(\picorv32_core/n358 [21]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [21]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b22  (
    .clk(clk),
    .d(\picorv32_core/n358 [22]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [22]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b23  (
    .clk(clk),
    .d(\picorv32_core/n358 [23]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [23]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b24  (
    .clk(clk),
    .d(\picorv32_core/n358 [24]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [24]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b25  (
    .clk(clk),
    .d(\picorv32_core/n358 [25]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [25]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b26  (
    .clk(clk),
    .d(\picorv32_core/n358 [26]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [26]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b27  (
    .clk(clk),
    .d(\picorv32_core/n358 [27]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [27]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b28  (
    .clk(clk),
    .d(\picorv32_core/n358 [28]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [28]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b29  (
    .clk(clk),
    .d(\picorv32_core/n358 [29]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [29]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b3  (
    .clk(clk),
    .d(\picorv32_core/n358 [3]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [3]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b30  (
    .clk(clk),
    .d(\picorv32_core/n358 [30]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [30]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b31  (
    .clk(clk),
    .d(\picorv32_core/n358 [31]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [31]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b4  (
    .clk(clk),
    .d(\picorv32_core/n358 [4]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [4]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b5  (
    .clk(clk),
    .d(\picorv32_core/n358 [5]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [5]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b6  (
    .clk(clk),
    .d(\picorv32_core/n358 [6]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [6]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b7  (
    .clk(clk),
    .d(\picorv32_core/n358 [7]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [7]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b8  (
    .clk(clk),
    .d(\picorv32_core/n358 [8]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [8]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg11_b9  (
    .clk(clk),
    .d(\picorv32_core/n358 [9]),
    .en(\picorv32_core/n274 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm [9]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg12_b0  (
    .clk(clk),
    .d(\picorv32_core/n726 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_sh [0]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg12_b1  (
    .clk(clk),
    .d(\picorv32_core/n726 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_sh [1]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg12_b2  (
    .clk(clk),
    .d(\picorv32_core/n726 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_sh [2]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg12_b3  (
    .clk(clk),
    .d(\picorv32_core/n726 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_sh [3]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg12_b4  (
    .clk(clk),
    .d(\picorv32_core/n726 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_sh [4]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b0  (
    .clk(clk),
    .d(\picorv32_core/n725 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [0]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b1  (
    .clk(clk),
    .d(\picorv32_core/n725 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [1]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b10  (
    .clk(clk),
    .d(\picorv32_core/n725 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [10]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b11  (
    .clk(clk),
    .d(\picorv32_core/n725 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [11]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b12  (
    .clk(clk),
    .d(\picorv32_core/n725 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [12]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b13  (
    .clk(clk),
    .d(\picorv32_core/n725 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [13]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b14  (
    .clk(clk),
    .d(\picorv32_core/n725 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [14]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b15  (
    .clk(clk),
    .d(\picorv32_core/n725 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [15]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b16  (
    .clk(clk),
    .d(\picorv32_core/n725 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [16]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b17  (
    .clk(clk),
    .d(\picorv32_core/n725 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [17]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b18  (
    .clk(clk),
    .d(\picorv32_core/n725 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [18]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b19  (
    .clk(clk),
    .d(\picorv32_core/n725 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [19]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b2  (
    .clk(clk),
    .d(\picorv32_core/n725 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [2]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b20  (
    .clk(clk),
    .d(\picorv32_core/n725 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [20]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b21  (
    .clk(clk),
    .d(\picorv32_core/n725 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [21]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b22  (
    .clk(clk),
    .d(\picorv32_core/n725 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [22]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b23  (
    .clk(clk),
    .d(\picorv32_core/n725 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [23]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b24  (
    .clk(clk),
    .d(\picorv32_core/n725 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [24]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b25  (
    .clk(clk),
    .d(\picorv32_core/n725 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [25]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b26  (
    .clk(clk),
    .d(\picorv32_core/n725 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [26]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b27  (
    .clk(clk),
    .d(\picorv32_core/n725 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [27]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b28  (
    .clk(clk),
    .d(\picorv32_core/n725 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [28]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b29  (
    .clk(clk),
    .d(\picorv32_core/n725 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [29]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b3  (
    .clk(clk),
    .d(\picorv32_core/n725 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [3]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b30  (
    .clk(clk),
    .d(\picorv32_core/n725 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [30]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b31  (
    .clk(clk),
    .d(\picorv32_core/n725 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [31]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b4  (
    .clk(clk),
    .d(\picorv32_core/n725 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [4]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b5  (
    .clk(clk),
    .d(\picorv32_core/n725 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [5]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b6  (
    .clk(clk),
    .d(\picorv32_core/n725 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [6]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b7  (
    .clk(clk),
    .d(\picorv32_core/n725 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [7]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b8  (
    .clk(clk),
    .d(\picorv32_core/n725 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [8]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg13_b9  (
    .clk(clk),
    .d(\picorv32_core/n725 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/reg_out [9]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b0  (
    .clk(clk),
    .d(\picorv32_core/alu_out [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [0]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b1  (
    .clk(clk),
    .d(\picorv32_core/alu_out [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [1]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b10  (
    .clk(clk),
    .d(\picorv32_core/alu_out [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [10]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b11  (
    .clk(clk),
    .d(\picorv32_core/alu_out [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [11]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b12  (
    .clk(clk),
    .d(\picorv32_core/alu_out [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [12]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b13  (
    .clk(clk),
    .d(\picorv32_core/alu_out [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [13]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b14  (
    .clk(clk),
    .d(\picorv32_core/alu_out [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [14]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b15  (
    .clk(clk),
    .d(\picorv32_core/alu_out [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [15]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b16  (
    .clk(clk),
    .d(\picorv32_core/alu_out [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [16]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b17  (
    .clk(clk),
    .d(\picorv32_core/alu_out [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [17]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b18  (
    .clk(clk),
    .d(\picorv32_core/alu_out [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [18]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b19  (
    .clk(clk),
    .d(\picorv32_core/alu_out [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [19]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b2  (
    .clk(clk),
    .d(\picorv32_core/alu_out [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [2]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b20  (
    .clk(clk),
    .d(\picorv32_core/alu_out [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [20]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b21  (
    .clk(clk),
    .d(\picorv32_core/alu_out [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [21]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b22  (
    .clk(clk),
    .d(\picorv32_core/alu_out [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [22]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b23  (
    .clk(clk),
    .d(\picorv32_core/alu_out [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [23]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b24  (
    .clk(clk),
    .d(\picorv32_core/alu_out [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [24]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b25  (
    .clk(clk),
    .d(\picorv32_core/alu_out [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [25]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b26  (
    .clk(clk),
    .d(\picorv32_core/alu_out [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [26]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b27  (
    .clk(clk),
    .d(\picorv32_core/alu_out [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [27]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b28  (
    .clk(clk),
    .d(\picorv32_core/alu_out [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [28]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b29  (
    .clk(clk),
    .d(\picorv32_core/alu_out [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [29]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b3  (
    .clk(clk),
    .d(\picorv32_core/alu_out [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [3]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b30  (
    .clk(clk),
    .d(\picorv32_core/alu_out [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [30]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b31  (
    .clk(clk),
    .d(\picorv32_core/alu_out [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [31]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b4  (
    .clk(clk),
    .d(\picorv32_core/alu_out [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [4]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b5  (
    .clk(clk),
    .d(\picorv32_core/alu_out [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [5]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b6  (
    .clk(clk),
    .d(\picorv32_core/alu_out [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [6]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b7  (
    .clk(clk),
    .d(\picorv32_core/alu_out [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [7]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b8  (
    .clk(clk),
    .d(\picorv32_core/alu_out [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [8]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg14_b9  (
    .clk(clk),
    .d(\picorv32_core/alu_out [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/alu_out_q [9]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b0  (
    .clk(clk),
    .d(\picorv32_core/n459 [0]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [0]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b1  (
    .clk(clk),
    .d(\picorv32_core/n459 [1]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [1]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b10  (
    .clk(clk),
    .d(\picorv32_core/n459 [10]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [10]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b11  (
    .clk(clk),
    .d(\picorv32_core/n459 [11]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [11]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b12  (
    .clk(clk),
    .d(\picorv32_core/n459 [12]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [12]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b13  (
    .clk(clk),
    .d(\picorv32_core/n459 [13]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [13]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b14  (
    .clk(clk),
    .d(\picorv32_core/n459 [14]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [14]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b15  (
    .clk(clk),
    .d(\picorv32_core/n459 [15]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [15]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b16  (
    .clk(clk),
    .d(\picorv32_core/n459 [16]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [16]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b17  (
    .clk(clk),
    .d(\picorv32_core/n459 [17]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [17]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b18  (
    .clk(clk),
    .d(\picorv32_core/n459 [18]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [18]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b19  (
    .clk(clk),
    .d(\picorv32_core/n459 [19]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [19]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b2  (
    .clk(clk),
    .d(\picorv32_core/n459 [2]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [2]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b20  (
    .clk(clk),
    .d(\picorv32_core/n459 [20]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [20]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b21  (
    .clk(clk),
    .d(\picorv32_core/n459 [21]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [21]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b22  (
    .clk(clk),
    .d(\picorv32_core/n459 [22]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [22]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b23  (
    .clk(clk),
    .d(\picorv32_core/n459 [23]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [23]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b24  (
    .clk(clk),
    .d(\picorv32_core/n459 [24]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [24]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b25  (
    .clk(clk),
    .d(\picorv32_core/n459 [25]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [25]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b26  (
    .clk(clk),
    .d(\picorv32_core/n459 [26]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [26]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b27  (
    .clk(clk),
    .d(\picorv32_core/n459 [27]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [27]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b28  (
    .clk(clk),
    .d(\picorv32_core/n459 [28]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [28]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b29  (
    .clk(clk),
    .d(\picorv32_core/n459 [29]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [29]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b3  (
    .clk(clk),
    .d(\picorv32_core/n459 [3]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [3]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b30  (
    .clk(clk),
    .d(\picorv32_core/n459 [30]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [30]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b31  (
    .clk(clk),
    .d(\picorv32_core/n459 [31]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [31]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b32  (
    .clk(clk),
    .d(\picorv32_core/n459 [32]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [32]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b33  (
    .clk(clk),
    .d(\picorv32_core/n459 [33]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [33]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b34  (
    .clk(clk),
    .d(\picorv32_core/n459 [34]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [34]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b35  (
    .clk(clk),
    .d(\picorv32_core/n459 [35]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [35]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b36  (
    .clk(clk),
    .d(\picorv32_core/n459 [36]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [36]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b37  (
    .clk(clk),
    .d(\picorv32_core/n459 [37]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [37]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b38  (
    .clk(clk),
    .d(\picorv32_core/n459 [38]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [38]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b39  (
    .clk(clk),
    .d(\picorv32_core/n459 [39]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [39]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b4  (
    .clk(clk),
    .d(\picorv32_core/n459 [4]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [4]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b40  (
    .clk(clk),
    .d(\picorv32_core/n459 [40]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [40]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b41  (
    .clk(clk),
    .d(\picorv32_core/n459 [41]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [41]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b42  (
    .clk(clk),
    .d(\picorv32_core/n459 [42]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [42]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b43  (
    .clk(clk),
    .d(\picorv32_core/n459 [43]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [43]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b44  (
    .clk(clk),
    .d(\picorv32_core/n459 [44]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [44]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b45  (
    .clk(clk),
    .d(\picorv32_core/n459 [45]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [45]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b46  (
    .clk(clk),
    .d(\picorv32_core/n459 [46]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [46]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b47  (
    .clk(clk),
    .d(\picorv32_core/n459 [47]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [47]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b48  (
    .clk(clk),
    .d(\picorv32_core/n459 [48]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [48]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b49  (
    .clk(clk),
    .d(\picorv32_core/n459 [49]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [49]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b5  (
    .clk(clk),
    .d(\picorv32_core/n459 [5]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [5]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b50  (
    .clk(clk),
    .d(\picorv32_core/n459 [50]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [50]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b51  (
    .clk(clk),
    .d(\picorv32_core/n459 [51]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [51]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b52  (
    .clk(clk),
    .d(\picorv32_core/n459 [52]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [52]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b53  (
    .clk(clk),
    .d(\picorv32_core/n459 [53]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [53]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b54  (
    .clk(clk),
    .d(\picorv32_core/n459 [54]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [54]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b55  (
    .clk(clk),
    .d(\picorv32_core/n459 [55]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [55]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b56  (
    .clk(clk),
    .d(\picorv32_core/n459 [56]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [56]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b57  (
    .clk(clk),
    .d(\picorv32_core/n459 [57]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [57]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b58  (
    .clk(clk),
    .d(\picorv32_core/n459 [58]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [58]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b59  (
    .clk(clk),
    .d(\picorv32_core/n459 [59]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [59]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b6  (
    .clk(clk),
    .d(\picorv32_core/n459 [6]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [6]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b60  (
    .clk(clk),
    .d(\picorv32_core/n459 [60]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [60]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b61  (
    .clk(clk),
    .d(\picorv32_core/n459 [61]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [61]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b62  (
    .clk(clk),
    .d(\picorv32_core/n459 [62]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [62]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b63  (
    .clk(clk),
    .d(\picorv32_core/n459 [63]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [63]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b7  (
    .clk(clk),
    .d(\picorv32_core/n459 [7]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [7]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b8  (
    .clk(clk),
    .d(\picorv32_core/n459 [8]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [8]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg15_b9  (
    .clk(clk),
    .d(\picorv32_core/n459 [9]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_cycle [9]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b0  (
    .clk(clk),
    .d(\picorv32_core/n500 [0]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [0]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b1  (
    .clk(clk),
    .d(\picorv32_core/n500 [1]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [1]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b10  (
    .clk(clk),
    .d(\picorv32_core/n500 [10]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [10]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b11  (
    .clk(clk),
    .d(\picorv32_core/n500 [11]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [11]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b12  (
    .clk(clk),
    .d(\picorv32_core/n500 [12]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [12]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b13  (
    .clk(clk),
    .d(\picorv32_core/n500 [13]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [13]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b14  (
    .clk(clk),
    .d(\picorv32_core/n500 [14]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [14]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b15  (
    .clk(clk),
    .d(\picorv32_core/n500 [15]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [15]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b16  (
    .clk(clk),
    .d(\picorv32_core/n500 [16]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [16]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b17  (
    .clk(clk),
    .d(\picorv32_core/n500 [17]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [17]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b18  (
    .clk(clk),
    .d(\picorv32_core/n500 [18]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [18]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b19  (
    .clk(clk),
    .d(\picorv32_core/n500 [19]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [19]));  // ../src/picorv32.v(1906)
  reg_ar_ss_w1 \picorv32_core/reg17_b2  (
    .clk(clk),
    .d(\picorv32_core/n500 [2]),
    .en(\picorv32_core/n663 ),
    .reset(1'b0),
    .set(~resetn),
    .q(\picorv32_core/reg_pc [2]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b20  (
    .clk(clk),
    .d(\picorv32_core/n500 [20]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [20]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b21  (
    .clk(clk),
    .d(\picorv32_core/n500 [21]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [21]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b22  (
    .clk(clk),
    .d(\picorv32_core/n500 [22]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [22]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b23  (
    .clk(clk),
    .d(\picorv32_core/n500 [23]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [23]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b24  (
    .clk(clk),
    .d(\picorv32_core/n500 [24]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [24]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b25  (
    .clk(clk),
    .d(\picorv32_core/n500 [25]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [25]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b26  (
    .clk(clk),
    .d(\picorv32_core/n500 [26]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [26]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b27  (
    .clk(clk),
    .d(\picorv32_core/n500 [27]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [27]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b28  (
    .clk(clk),
    .d(\picorv32_core/n500 [28]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [28]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b29  (
    .clk(clk),
    .d(\picorv32_core/n500 [29]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [29]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b3  (
    .clk(clk),
    .d(\picorv32_core/n500 [3]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [3]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b30  (
    .clk(clk),
    .d(\picorv32_core/n500 [30]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [30]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b31  (
    .clk(clk),
    .d(\picorv32_core/n500 [31]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [31]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b4  (
    .clk(clk),
    .d(\picorv32_core/n500 [4]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [4]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b5  (
    .clk(clk),
    .d(\picorv32_core/n500 [5]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [5]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b6  (
    .clk(clk),
    .d(\picorv32_core/n500 [6]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [6]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b7  (
    .clk(clk),
    .d(\picorv32_core/n500 [7]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [7]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b8  (
    .clk(clk),
    .d(\picorv32_core/n500 [8]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [8]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg17_b9  (
    .clk(clk),
    .d(\picorv32_core/n500 [9]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_pc [9]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b0  (
    .clk(clk),
    .d(\picorv32_core/n511 [0]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [0]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b1  (
    .clk(clk),
    .d(\picorv32_core/n511 [1]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [1]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b10  (
    .clk(clk),
    .d(\picorv32_core/n511 [10]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [10]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b11  (
    .clk(clk),
    .d(\picorv32_core/n511 [11]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [11]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b12  (
    .clk(clk),
    .d(\picorv32_core/n511 [12]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [12]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b13  (
    .clk(clk),
    .d(\picorv32_core/n511 [13]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [13]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b14  (
    .clk(clk),
    .d(\picorv32_core/n511 [14]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [14]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b15  (
    .clk(clk),
    .d(\picorv32_core/n511 [15]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [15]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b16  (
    .clk(clk),
    .d(\picorv32_core/n511 [16]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [16]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b17  (
    .clk(clk),
    .d(\picorv32_core/n511 [17]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [17]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b18  (
    .clk(clk),
    .d(\picorv32_core/n511 [18]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [18]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b19  (
    .clk(clk),
    .d(\picorv32_core/n511 [19]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [19]));  // ../src/picorv32.v(1906)
  reg_ar_ss_w1 \picorv32_core/reg18_b2  (
    .clk(clk),
    .d(\picorv32_core/n511 [2]),
    .en(\picorv32_core/n663 ),
    .reset(1'b0),
    .set(~resetn),
    .q(\picorv32_core/reg_next_pc [2]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b20  (
    .clk(clk),
    .d(\picorv32_core/n511 [20]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [20]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b21  (
    .clk(clk),
    .d(\picorv32_core/n511 [21]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [21]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b22  (
    .clk(clk),
    .d(\picorv32_core/n511 [22]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [22]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b23  (
    .clk(clk),
    .d(\picorv32_core/n511 [23]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [23]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b24  (
    .clk(clk),
    .d(\picorv32_core/n511 [24]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [24]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b25  (
    .clk(clk),
    .d(\picorv32_core/n511 [25]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [25]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b26  (
    .clk(clk),
    .d(\picorv32_core/n511 [26]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [26]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b27  (
    .clk(clk),
    .d(\picorv32_core/n511 [27]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [27]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b28  (
    .clk(clk),
    .d(\picorv32_core/n511 [28]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [28]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b29  (
    .clk(clk),
    .d(\picorv32_core/n511 [29]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [29]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b3  (
    .clk(clk),
    .d(\picorv32_core/n511 [3]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [3]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b30  (
    .clk(clk),
    .d(\picorv32_core/n511 [30]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [30]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b31  (
    .clk(clk),
    .d(\picorv32_core/n511 [31]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [31]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b4  (
    .clk(clk),
    .d(\picorv32_core/n511 [4]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [4]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b5  (
    .clk(clk),
    .d(\picorv32_core/n511 [5]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [5]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b6  (
    .clk(clk),
    .d(\picorv32_core/n511 [6]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [6]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b7  (
    .clk(clk),
    .d(\picorv32_core/n511 [7]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [7]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b8  (
    .clk(clk),
    .d(\picorv32_core/n511 [8]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [8]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg18_b9  (
    .clk(clk),
    .d(\picorv32_core/n511 [9]),
    .en(\picorv32_core/n663 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/reg_next_pc [9]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b0  (
    .clk(clk),
    .d(\picorv32_core/n503 [0]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [0]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b1  (
    .clk(clk),
    .d(\picorv32_core/n503 [1]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [1]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b10  (
    .clk(clk),
    .d(\picorv32_core/n503 [10]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [10]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b11  (
    .clk(clk),
    .d(\picorv32_core/n503 [11]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [11]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b12  (
    .clk(clk),
    .d(\picorv32_core/n503 [12]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [12]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b13  (
    .clk(clk),
    .d(\picorv32_core/n503 [13]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [13]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b14  (
    .clk(clk),
    .d(\picorv32_core/n503 [14]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [14]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b15  (
    .clk(clk),
    .d(\picorv32_core/n503 [15]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [15]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b16  (
    .clk(clk),
    .d(\picorv32_core/n503 [16]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [16]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b17  (
    .clk(clk),
    .d(\picorv32_core/n503 [17]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [17]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b18  (
    .clk(clk),
    .d(\picorv32_core/n503 [18]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [18]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b19  (
    .clk(clk),
    .d(\picorv32_core/n503 [19]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [19]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b2  (
    .clk(clk),
    .d(\picorv32_core/n503 [2]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [2]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b20  (
    .clk(clk),
    .d(\picorv32_core/n503 [20]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [20]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b21  (
    .clk(clk),
    .d(\picorv32_core/n503 [21]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [21]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b22  (
    .clk(clk),
    .d(\picorv32_core/n503 [22]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [22]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b23  (
    .clk(clk),
    .d(\picorv32_core/n503 [23]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [23]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b24  (
    .clk(clk),
    .d(\picorv32_core/n503 [24]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [24]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b25  (
    .clk(clk),
    .d(\picorv32_core/n503 [25]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [25]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b26  (
    .clk(clk),
    .d(\picorv32_core/n503 [26]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [26]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b27  (
    .clk(clk),
    .d(\picorv32_core/n503 [27]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [27]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b28  (
    .clk(clk),
    .d(\picorv32_core/n503 [28]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [28]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b29  (
    .clk(clk),
    .d(\picorv32_core/n503 [29]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [29]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b3  (
    .clk(clk),
    .d(\picorv32_core/n503 [3]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [3]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b30  (
    .clk(clk),
    .d(\picorv32_core/n503 [30]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [30]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b31  (
    .clk(clk),
    .d(\picorv32_core/n503 [31]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [31]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b32  (
    .clk(clk),
    .d(\picorv32_core/n503 [32]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [32]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b33  (
    .clk(clk),
    .d(\picorv32_core/n503 [33]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [33]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b34  (
    .clk(clk),
    .d(\picorv32_core/n503 [34]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [34]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b35  (
    .clk(clk),
    .d(\picorv32_core/n503 [35]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [35]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b36  (
    .clk(clk),
    .d(\picorv32_core/n503 [36]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [36]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b37  (
    .clk(clk),
    .d(\picorv32_core/n503 [37]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [37]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b38  (
    .clk(clk),
    .d(\picorv32_core/n503 [38]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [38]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b39  (
    .clk(clk),
    .d(\picorv32_core/n503 [39]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [39]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b4  (
    .clk(clk),
    .d(\picorv32_core/n503 [4]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [4]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b40  (
    .clk(clk),
    .d(\picorv32_core/n503 [40]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [40]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b41  (
    .clk(clk),
    .d(\picorv32_core/n503 [41]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [41]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b42  (
    .clk(clk),
    .d(\picorv32_core/n503 [42]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [42]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b43  (
    .clk(clk),
    .d(\picorv32_core/n503 [43]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [43]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b44  (
    .clk(clk),
    .d(\picorv32_core/n503 [44]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [44]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b45  (
    .clk(clk),
    .d(\picorv32_core/n503 [45]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [45]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b46  (
    .clk(clk),
    .d(\picorv32_core/n503 [46]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [46]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b47  (
    .clk(clk),
    .d(\picorv32_core/n503 [47]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [47]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b48  (
    .clk(clk),
    .d(\picorv32_core/n503 [48]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [48]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b49  (
    .clk(clk),
    .d(\picorv32_core/n503 [49]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [49]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b5  (
    .clk(clk),
    .d(\picorv32_core/n503 [5]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [5]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b50  (
    .clk(clk),
    .d(\picorv32_core/n503 [50]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [50]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b51  (
    .clk(clk),
    .d(\picorv32_core/n503 [51]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [51]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b52  (
    .clk(clk),
    .d(\picorv32_core/n503 [52]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [52]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b53  (
    .clk(clk),
    .d(\picorv32_core/n503 [53]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [53]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b54  (
    .clk(clk),
    .d(\picorv32_core/n503 [54]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [54]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b55  (
    .clk(clk),
    .d(\picorv32_core/n503 [55]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [55]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b56  (
    .clk(clk),
    .d(\picorv32_core/n503 [56]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [56]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b57  (
    .clk(clk),
    .d(\picorv32_core/n503 [57]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [57]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b58  (
    .clk(clk),
    .d(\picorv32_core/n503 [58]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [58]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b59  (
    .clk(clk),
    .d(\picorv32_core/n503 [59]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [59]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b6  (
    .clk(clk),
    .d(\picorv32_core/n503 [6]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [6]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b60  (
    .clk(clk),
    .d(\picorv32_core/n503 [60]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [60]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b61  (
    .clk(clk),
    .d(\picorv32_core/n503 [61]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [61]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b62  (
    .clk(clk),
    .d(\picorv32_core/n503 [62]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [62]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b63  (
    .clk(clk),
    .d(\picorv32_core/n503 [63]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [63]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b7  (
    .clk(clk),
    .d(\picorv32_core/n503 [7]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [7]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b8  (
    .clk(clk),
    .d(\picorv32_core/n503 [8]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [8]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg19_b9  (
    .clk(clk),
    .d(\picorv32_core/n503 [9]),
    .en(\picorv32_core/sel39_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\picorv32_core/count_instr [9]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg1_b0  (
    .clk(clk),
    .d(\picorv32_core/n154 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_state [0]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg1_b1  (
    .clk(clk),
    .d(\picorv32_core/n154 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_state [1]));  // ../src/picorv32.v(605)
  reg_sr_as_w1 \picorv32_core/reg22_b0  (
    .clk(clk),
    .d(\picorv32_core/n716 [0]),
    .en(1'b1),
    .reset(~\picorv32_core/mux164_b0_sel_is_0_o ),
    .set(1'b0),
    .q(\picorv32_core/cpu_state [0]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg22_b1  (
    .clk(clk),
    .d(\picorv32_core/n716 [1]),
    .en(1'b1),
    .reset(~\picorv32_core/mux164_b0_sel_is_0_o ),
    .set(1'b0),
    .q(\picorv32_core/cpu_state [1]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg22_b2  (
    .clk(clk),
    .d(\picorv32_core/n716 [2]),
    .en(1'b1),
    .reset(~\picorv32_core/mux164_b0_sel_is_0_o ),
    .set(1'b0),
    .q(\picorv32_core/cpu_state [2]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg22_b3  (
    .clk(clk),
    .d(\picorv32_core/n716 [3]),
    .en(1'b1),
    .reset(~\picorv32_core/mux164_b0_sel_is_0_o ),
    .set(1'b0),
    .q(\picorv32_core/cpu_state [3]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg22_b4  (
    .clk(clk),
    .d(\picorv32_core/n716 [4]),
    .en(1'b1),
    .reset(~\picorv32_core/mux164_b0_sel_is_0_o ),
    .set(1'b0),
    .q(\picorv32_core/cpu_state [4]));  // ../src/picorv32.v(1906)
  reg_sr_as_w1 \picorv32_core/reg22_b5  (
    .clk(clk),
    .d(\picorv32_core/n716 [5]),
    .en(1'b1),
    .reset(~\picorv32_core/mux164_b0_sel_is_0_o ),
    .set(1'b0),
    .q(\picorv32_core/cpu_state [5]));  // ../src/picorv32.v(1906)
  reg_sr_ss_w1 \picorv32_core/reg22_b6  (
    .clk(clk),
    .d(\picorv32_core/n692 [6]),
    .en(1'b1),
    .reset(~\picorv32_core/mux164_b0_sel_is_0_o ),
    .set(~resetn),
    .q(\picorv32_core/cpu_state [6]));  // ../src/picorv32.v(1906)
  reg_ar_ss_w1 \picorv32_core/reg22_b7  (
    .clk(clk),
    .d(\picorv32_core/n716 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(~\picorv32_core/mux164_b0_sel_is_0_o ),
    .q(\picorv32_core/cpu_state [7]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg23_b0  (
    .clk(clk),
    .d(\picorv32_core/n672 [0]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_wordsize [0]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg23_b1  (
    .clk(clk),
    .d(\picorv32_core/n672 [1]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_wordsize [1]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg24_b0  (
    .clk(clk),
    .d(\picorv32_core/n688 [0]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/latched_rd [0]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg24_b1  (
    .clk(clk),
    .d(\picorv32_core/n688 [1]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/latched_rd [1]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg24_b2  (
    .clk(clk),
    .d(\picorv32_core/n688 [2]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/latched_rd [2]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg24_b3  (
    .clk(clk),
    .d(\picorv32_core/n688 [3]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/latched_rd [3]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg24_b4  (
    .clk(clk),
    .d(\picorv32_core/n688 [4]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/latched_rd [4]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b0  (
    .clk(clk),
    .d(\picorv32_core/n693 [0]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$0$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b1  (
    .clk(clk),
    .d(\picorv32_core/n693 [1]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$1$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b10  (
    .clk(clk),
    .d(\picorv32_core/n693 [10]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$10$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b11  (
    .clk(clk),
    .d(\picorv32_core/n693 [11]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$11$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b12  (
    .clk(clk),
    .d(\picorv32_core/n693 [12]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$12$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b13  (
    .clk(clk),
    .d(\picorv32_core/n693 [13]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$13$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b14  (
    .clk(clk),
    .d(\picorv32_core/n693 [14]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$14$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b15  (
    .clk(clk),
    .d(\picorv32_core/n693 [15]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$15$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b16  (
    .clk(clk),
    .d(\picorv32_core/n693 [16]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$16$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b17  (
    .clk(clk),
    .d(\picorv32_core/n693 [17]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$17$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b18  (
    .clk(clk),
    .d(\picorv32_core/n693 [18]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$18$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b19  (
    .clk(clk),
    .d(\picorv32_core/n693 [19]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$19$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b2  (
    .clk(clk),
    .d(\picorv32_core/n693 [2]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$2$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b20  (
    .clk(clk),
    .d(\picorv32_core/n693 [20]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$20$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b21  (
    .clk(clk),
    .d(\picorv32_core/n693 [21]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$21$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b22  (
    .clk(clk),
    .d(\picorv32_core/n693 [22]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$22$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b23  (
    .clk(clk),
    .d(\picorv32_core/n693 [23]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$23$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b24  (
    .clk(clk),
    .d(\picorv32_core/n693 [24]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$24$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b25  (
    .clk(clk),
    .d(\picorv32_core/n693 [25]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$25$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b26  (
    .clk(clk),
    .d(\picorv32_core/n693 [26]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$26$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b27  (
    .clk(clk),
    .d(\picorv32_core/n693 [27]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$27$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b28  (
    .clk(clk),
    .d(\picorv32_core/n693 [28]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$28$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b29  (
    .clk(clk),
    .d(\picorv32_core/n693 [29]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$29$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b3  (
    .clk(clk),
    .d(\picorv32_core/n693 [3]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$3$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b30  (
    .clk(clk),
    .d(\picorv32_core/n693 [30]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$30$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b31  (
    .clk(clk),
    .d(\picorv32_core/n693 [31]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$31$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b4  (
    .clk(clk),
    .d(\picorv32_core/n693 [4]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$4$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b5  (
    .clk(clk),
    .d(\picorv32_core/n693 [5]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$5$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b6  (
    .clk(clk),
    .d(\picorv32_core/n693 [6]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$6$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b7  (
    .clk(clk),
    .d(\picorv32_core/n693 [7]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$7$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b8  (
    .clk(clk),
    .d(\picorv32_core/n693 [8]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$8$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg25_b9  (
    .clk(clk),
    .d(\picorv32_core/n693 [9]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs1$9$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b0  (
    .clk(clk),
    .d(\picorv32_core/n694 [0]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(mem_la_wdata[0]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b1  (
    .clk(clk),
    .d(\picorv32_core/n694 [1]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(mem_la_wdata[1]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b10  (
    .clk(clk),
    .d(\picorv32_core/n694 [10]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$10$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b11  (
    .clk(clk),
    .d(\picorv32_core/n694 [11]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$11$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b12  (
    .clk(clk),
    .d(\picorv32_core/n694 [12]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$12$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b13  (
    .clk(clk),
    .d(\picorv32_core/n694 [13]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$13$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b14  (
    .clk(clk),
    .d(\picorv32_core/n694 [14]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$14$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b15  (
    .clk(clk),
    .d(\picorv32_core/n694 [15]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$15$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b16  (
    .clk(clk),
    .d(\picorv32_core/n694 [16]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$16$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b17  (
    .clk(clk),
    .d(\picorv32_core/n694 [17]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$17$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b18  (
    .clk(clk),
    .d(\picorv32_core/n694 [18]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$18$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b19  (
    .clk(clk),
    .d(\picorv32_core/n694 [19]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$19$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b2  (
    .clk(clk),
    .d(\picorv32_core/n694 [2]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(mem_la_wdata[2]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b20  (
    .clk(clk),
    .d(\picorv32_core/n694 [20]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$20$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b21  (
    .clk(clk),
    .d(\picorv32_core/n694 [21]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$21$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b22  (
    .clk(clk),
    .d(\picorv32_core/n694 [22]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$22$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b23  (
    .clk(clk),
    .d(\picorv32_core/n694 [23]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$23$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b24  (
    .clk(clk),
    .d(\picorv32_core/n694 [24]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$24$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b25  (
    .clk(clk),
    .d(\picorv32_core/n694 [25]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$25$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b26  (
    .clk(clk),
    .d(\picorv32_core/n694 [26]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$26$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b27  (
    .clk(clk),
    .d(\picorv32_core/n694 [27]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$27$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b28  (
    .clk(clk),
    .d(\picorv32_core/n694 [28]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$28$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b29  (
    .clk(clk),
    .d(\picorv32_core/n694 [29]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$29$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b3  (
    .clk(clk),
    .d(\picorv32_core/n694 [3]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(mem_la_wdata[3]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b30  (
    .clk(clk),
    .d(\picorv32_core/n694 [30]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$30$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b31  (
    .clk(clk),
    .d(\picorv32_core/n694 [31]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$31$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b4  (
    .clk(clk),
    .d(\picorv32_core/n694 [4]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(mem_la_wdata[4]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b5  (
    .clk(clk),
    .d(\picorv32_core/n694 [5]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(mem_la_wdata[5]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b6  (
    .clk(clk),
    .d(\picorv32_core/n694 [6]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(mem_la_wdata[6]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b7  (
    .clk(clk),
    .d(\picorv32_core/n694 [7]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(mem_la_wdata[7]));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b8  (
    .clk(clk),
    .d(\picorv32_core/n694 [8]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$8$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg26_b9  (
    .clk(clk),
    .d(\picorv32_core/n694 [9]),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/pcpi_rs2$9$ ));  // ../src/picorv32.v(1906)
  reg_ar_as_w1 \picorv32_core/reg5_b0  (
    .clk(clk),
    .d(\picorv32_core/n136 [0]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [0]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b1  (
    .clk(clk),
    .d(\picorv32_core/n136 [1]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [1]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b10  (
    .clk(clk),
    .d(\picorv32_core/n136 [10]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [10]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b11  (
    .clk(clk),
    .d(\picorv32_core/n136 [11]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [11]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b12  (
    .clk(clk),
    .d(\picorv32_core/n136 [12]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [12]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b13  (
    .clk(clk),
    .d(\picorv32_core/n136 [13]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [13]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b14  (
    .clk(clk),
    .d(\picorv32_core/n136 [14]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [14]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b15  (
    .clk(clk),
    .d(\picorv32_core/n136 [15]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [15]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b2  (
    .clk(clk),
    .d(\picorv32_core/n136 [2]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [2]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b3  (
    .clk(clk),
    .d(\picorv32_core/n136 [3]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [3]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b4  (
    .clk(clk),
    .d(\picorv32_core/n136 [4]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [4]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b5  (
    .clk(clk),
    .d(\picorv32_core/n136 [5]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [5]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b6  (
    .clk(clk),
    .d(\picorv32_core/n136 [6]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [6]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b7  (
    .clk(clk),
    .d(\picorv32_core/n136 [7]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [7]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b8  (
    .clk(clk),
    .d(\picorv32_core/n136 [8]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [8]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg5_b9  (
    .clk(clk),
    .d(\picorv32_core/n136 [9]),
    .en(\picorv32_core/mux68_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/mem_16bit_buffer [9]));  // ../src/picorv32.v(605)
  reg_ar_as_w1 \picorv32_core/reg6_b1  (
    .clk(clk),
    .d(\picorv32_core/n248 [0]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [1]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b10  (
    .clk(clk),
    .d(\picorv32_core/n248 [9]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [10]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b11  (
    .clk(clk),
    .d(\picorv32_core/n248 [10]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [11]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b12  (
    .clk(clk),
    .d(\picorv32_core/mem_rdata_latched [12]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [12]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b13  (
    .clk(clk),
    .d(\picorv32_core/n248 [11]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [13]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b14  (
    .clk(clk),
    .d(\picorv32_core/n248 [12]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [14]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b15  (
    .clk(clk),
    .d(\picorv32_core/n248 [13]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [15]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b16  (
    .clk(clk),
    .d(\picorv32_core/n248 [14]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [16]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b17  (
    .clk(clk),
    .d(\picorv32_core/n248 [15]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [17]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b18  (
    .clk(clk),
    .d(\picorv32_core/n248 [16]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [18]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b19  (
    .clk(clk),
    .d(\picorv32_core/n248 [17]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [19]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b2  (
    .clk(clk),
    .d(\picorv32_core/n248 [1]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [2]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b20  (
    .clk(clk),
    .d(\picorv32_core/n248 [18]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [20]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b3  (
    .clk(clk),
    .d(\picorv32_core/n248 [2]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [3]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b4  (
    .clk(clk),
    .d(\picorv32_core/n248 [3]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [4]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b5  (
    .clk(clk),
    .d(\picorv32_core/n248 [4]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [5]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b6  (
    .clk(clk),
    .d(\picorv32_core/n248 [5]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [6]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b7  (
    .clk(clk),
    .d(\picorv32_core/n248 [6]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [7]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b8  (
    .clk(clk),
    .d(\picorv32_core/n248 [7]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [8]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg6_b9  (
    .clk(clk),
    .d(\picorv32_core/n248 [8]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_imm_uj [9]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg7_b0  (
    .clk(clk),
    .d(\picorv32_core/n245 [0]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rd [0]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg7_b1  (
    .clk(clk),
    .d(\picorv32_core/n245 [1]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rd [1]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg7_b2  (
    .clk(clk),
    .d(\picorv32_core/n245 [2]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rd [2]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg7_b3  (
    .clk(clk),
    .d(\picorv32_core/n245 [3]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rd [3]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg7_b4  (
    .clk(clk),
    .d(\picorv32_core/n245 [4]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rd [4]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg8_b0  (
    .clk(clk),
    .d(\picorv32_core/n246 [0]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rs1 [0]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg8_b1  (
    .clk(clk),
    .d(\picorv32_core/n246 [1]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rs1 [1]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg8_b2  (
    .clk(clk),
    .d(\picorv32_core/n246 [2]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rs1 [2]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg8_b3  (
    .clk(clk),
    .d(\picorv32_core/n246 [3]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rs1 [3]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg8_b4  (
    .clk(clk),
    .d(\picorv32_core/n246 [4]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rs1 [4]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg9_b0  (
    .clk(clk),
    .d(\picorv32_core/n247 [0]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rs2 [0]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg9_b1  (
    .clk(clk),
    .d(\picorv32_core/n247 [1]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rs2 [1]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg9_b2  (
    .clk(clk),
    .d(\picorv32_core/n247 [2]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rs2 [2]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg9_b3  (
    .clk(clk),
    .d(\picorv32_core/n247 [3]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rs2 [3]));  // ../src/picorv32.v(1120)
  reg_ar_as_w1 \picorv32_core/reg9_b4  (
    .clk(clk),
    .d(\picorv32_core/n247 [4]),
    .en(\picorv32_core/n170 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\picorv32_core/decoded_rs2 [4]));  // ../src/picorv32.v(1120)
  AL_MUX \picorv32_core/sel0_b0  (
    .i0(\picorv32_core/pcpi_rs1$4$ ),
    .i1(1'b0),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [0]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b1  (
    .i0(\picorv32_core/pcpi_rs1$5$ ),
    .i1(1'b0),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [1]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b10  (
    .i0(\picorv32_core/pcpi_rs1$14$ ),
    .i1(\picorv32_core/pcpi_rs1$6$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [10]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b11  (
    .i0(\picorv32_core/pcpi_rs1$15$ ),
    .i1(\picorv32_core/pcpi_rs1$7$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [11]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b12  (
    .i0(\picorv32_core/pcpi_rs1$16$ ),
    .i1(\picorv32_core/pcpi_rs1$8$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [12]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b13  (
    .i0(\picorv32_core/pcpi_rs1$17$ ),
    .i1(\picorv32_core/pcpi_rs1$9$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [13]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b14  (
    .i0(\picorv32_core/pcpi_rs1$18$ ),
    .i1(\picorv32_core/pcpi_rs1$10$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [14]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b15  (
    .i0(\picorv32_core/pcpi_rs1$19$ ),
    .i1(\picorv32_core/pcpi_rs1$11$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [15]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b16  (
    .i0(\picorv32_core/pcpi_rs1$20$ ),
    .i1(\picorv32_core/pcpi_rs1$12$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [16]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b17  (
    .i0(\picorv32_core/pcpi_rs1$21$ ),
    .i1(\picorv32_core/pcpi_rs1$13$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [17]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b18  (
    .i0(\picorv32_core/pcpi_rs1$22$ ),
    .i1(\picorv32_core/pcpi_rs1$14$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [18]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b19  (
    .i0(\picorv32_core/pcpi_rs1$23$ ),
    .i1(\picorv32_core/pcpi_rs1$15$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [19]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b2  (
    .i0(\picorv32_core/pcpi_rs1$6$ ),
    .i1(1'b0),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [2]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b20  (
    .i0(\picorv32_core/pcpi_rs1$24$ ),
    .i1(\picorv32_core/pcpi_rs1$16$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [20]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b21  (
    .i0(\picorv32_core/pcpi_rs1$25$ ),
    .i1(\picorv32_core/pcpi_rs1$17$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [21]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b22  (
    .i0(\picorv32_core/pcpi_rs1$26$ ),
    .i1(\picorv32_core/pcpi_rs1$18$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [22]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b23  (
    .i0(\picorv32_core/pcpi_rs1$27$ ),
    .i1(\picorv32_core/pcpi_rs1$19$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [23]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b24  (
    .i0(\picorv32_core/pcpi_rs1$28$ ),
    .i1(\picorv32_core/pcpi_rs1$20$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [24]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b25  (
    .i0(\picorv32_core/pcpi_rs1$29$ ),
    .i1(\picorv32_core/pcpi_rs1$21$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [25]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b26  (
    .i0(\picorv32_core/pcpi_rs1$30$ ),
    .i1(\picorv32_core/pcpi_rs1$22$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [26]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b27  (
    .i0(\picorv32_core/pcpi_rs1$31$ ),
    .i1(\picorv32_core/pcpi_rs1$23$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [27]));  // ../src/picorv32.v(1787)
  and \picorv32_core/sel0_b28/and_b0_0  (\picorv32_core/sel0_b28/B0 , \picorv32_core/pcpi_rs1$31$ , \picorv32_core/n557 );
  and \picorv32_core/sel0_b28/and_b0_2  (\picorv32_core/sel0_b28/B2 , \picorv32_core/pcpi_rs1$24$ , \picorv32_core/n555 );
  or \picorv32_core/sel0_b28/or_B0_or_B1_B2_o  (\picorv32_core/n558 [28], \picorv32_core/sel0_b28/B0 , \picorv32_core/sel0_b28/B2 );
  and \picorv32_core/sel0_b29/and_b0_2  (\picorv32_core/sel0_b29/B2 , \picorv32_core/pcpi_rs1$25$ , \picorv32_core/n555 );
  or \picorv32_core/sel0_b29/or_B0_or_B1_B2_o  (\picorv32_core/n558 [29], \picorv32_core/sel0_b28/B0 , \picorv32_core/sel0_b29/B2 );
  AL_MUX \picorv32_core/sel0_b3  (
    .i0(\picorv32_core/pcpi_rs1$7$ ),
    .i1(1'b0),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [3]));  // ../src/picorv32.v(1787)
  and \picorv32_core/sel0_b30/and_b0_2  (\picorv32_core/sel0_b30/B2 , \picorv32_core/pcpi_rs1$26$ , \picorv32_core/n555 );
  or \picorv32_core/sel0_b30/or_B0_or_B1_B2_o  (\picorv32_core/n558 [30], \picorv32_core/sel0_b28/B0 , \picorv32_core/sel0_b30/B2 );
  and \picorv32_core/sel0_b31/and_b0_2  (\picorv32_core/sel0_b31/B2 , \picorv32_core/pcpi_rs1$27$ , \picorv32_core/n555 );
  or \picorv32_core/sel0_b31/or_B0_or_B1_B2_o  (\picorv32_core/n558 [31], \picorv32_core/sel0_b28/B0 , \picorv32_core/sel0_b31/B2 );
  AL_MUX \picorv32_core/sel0_b32  (
    .i0(\picorv32_core/pcpi_rs1$1$ ),
    .i1(1'b0),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [0]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b33  (
    .i0(\picorv32_core/pcpi_rs1$2$ ),
    .i1(\picorv32_core/pcpi_rs1$0$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [1]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b34  (
    .i0(\picorv32_core/pcpi_rs1$3$ ),
    .i1(\picorv32_core/pcpi_rs1$1$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [2]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b35  (
    .i0(\picorv32_core/pcpi_rs1$4$ ),
    .i1(\picorv32_core/pcpi_rs1$2$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [3]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b36  (
    .i0(\picorv32_core/pcpi_rs1$5$ ),
    .i1(\picorv32_core/pcpi_rs1$3$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [4]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b37  (
    .i0(\picorv32_core/pcpi_rs1$6$ ),
    .i1(\picorv32_core/pcpi_rs1$4$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [5]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b38  (
    .i0(\picorv32_core/pcpi_rs1$7$ ),
    .i1(\picorv32_core/pcpi_rs1$5$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [6]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b39  (
    .i0(\picorv32_core/pcpi_rs1$8$ ),
    .i1(\picorv32_core/pcpi_rs1$6$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [7]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b4  (
    .i0(\picorv32_core/pcpi_rs1$8$ ),
    .i1(\picorv32_core/pcpi_rs1$0$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [4]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b40  (
    .i0(\picorv32_core/pcpi_rs1$9$ ),
    .i1(\picorv32_core/pcpi_rs1$7$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [8]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b41  (
    .i0(\picorv32_core/pcpi_rs1$10$ ),
    .i1(\picorv32_core/pcpi_rs1$8$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [9]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b42  (
    .i0(\picorv32_core/pcpi_rs1$11$ ),
    .i1(\picorv32_core/pcpi_rs1$9$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [10]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b43  (
    .i0(\picorv32_core/pcpi_rs1$12$ ),
    .i1(\picorv32_core/pcpi_rs1$10$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [11]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b44  (
    .i0(\picorv32_core/pcpi_rs1$13$ ),
    .i1(\picorv32_core/pcpi_rs1$11$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [12]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b45  (
    .i0(\picorv32_core/pcpi_rs1$14$ ),
    .i1(\picorv32_core/pcpi_rs1$12$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [13]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b46  (
    .i0(\picorv32_core/pcpi_rs1$15$ ),
    .i1(\picorv32_core/pcpi_rs1$13$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [14]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b47  (
    .i0(\picorv32_core/pcpi_rs1$16$ ),
    .i1(\picorv32_core/pcpi_rs1$14$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [15]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b48  (
    .i0(\picorv32_core/pcpi_rs1$17$ ),
    .i1(\picorv32_core/pcpi_rs1$15$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [16]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b49  (
    .i0(\picorv32_core/pcpi_rs1$18$ ),
    .i1(\picorv32_core/pcpi_rs1$16$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [17]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b5  (
    .i0(\picorv32_core/pcpi_rs1$9$ ),
    .i1(\picorv32_core/pcpi_rs1$1$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [5]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b50  (
    .i0(\picorv32_core/pcpi_rs1$19$ ),
    .i1(\picorv32_core/pcpi_rs1$17$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [18]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b51  (
    .i0(\picorv32_core/pcpi_rs1$20$ ),
    .i1(\picorv32_core/pcpi_rs1$18$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [19]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b52  (
    .i0(\picorv32_core/pcpi_rs1$21$ ),
    .i1(\picorv32_core/pcpi_rs1$19$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [20]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b53  (
    .i0(\picorv32_core/pcpi_rs1$22$ ),
    .i1(\picorv32_core/pcpi_rs1$20$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [21]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b54  (
    .i0(\picorv32_core/pcpi_rs1$23$ ),
    .i1(\picorv32_core/pcpi_rs1$21$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [22]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b55  (
    .i0(\picorv32_core/pcpi_rs1$24$ ),
    .i1(\picorv32_core/pcpi_rs1$22$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [23]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b56  (
    .i0(\picorv32_core/pcpi_rs1$25$ ),
    .i1(\picorv32_core/pcpi_rs1$23$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [24]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b57  (
    .i0(\picorv32_core/pcpi_rs1$26$ ),
    .i1(\picorv32_core/pcpi_rs1$24$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [25]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b58  (
    .i0(\picorv32_core/pcpi_rs1$27$ ),
    .i1(\picorv32_core/pcpi_rs1$25$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [26]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b59  (
    .i0(\picorv32_core/pcpi_rs1$28$ ),
    .i1(\picorv32_core/pcpi_rs1$26$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [27]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b6  (
    .i0(\picorv32_core/pcpi_rs1$10$ ),
    .i1(\picorv32_core/pcpi_rs1$2$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [6]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b60  (
    .i0(\picorv32_core/pcpi_rs1$29$ ),
    .i1(\picorv32_core/pcpi_rs1$27$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [28]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b61  (
    .i0(\picorv32_core/pcpi_rs1$30$ ),
    .i1(\picorv32_core/pcpi_rs1$28$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [29]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b62  (
    .i0(\picorv32_core/pcpi_rs1$31$ ),
    .i1(\picorv32_core/pcpi_rs1$29$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n563 [30]));  // ../src/picorv32.v(1787)
  and \picorv32_core/sel0_b63/and_b0_2  (\picorv32_core/sel0_b63/B2 , \picorv32_core/pcpi_rs1$30$ , \picorv32_core/n555 );
  or \picorv32_core/sel0_b63/or_B0_or_B1_B2_o  (\picorv32_core/n563 [31], \picorv32_core/sel0_b28/B0 , \picorv32_core/sel0_b63/B2 );
  AL_MUX \picorv32_core/sel0_b7  (
    .i0(\picorv32_core/pcpi_rs1$11$ ),
    .i1(\picorv32_core/pcpi_rs1$3$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [7]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b8  (
    .i0(\picorv32_core/pcpi_rs1$12$ ),
    .i1(\picorv32_core/pcpi_rs1$4$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [8]));  // ../src/picorv32.v(1787)
  AL_MUX \picorv32_core/sel0_b9  (
    .i0(\picorv32_core/pcpi_rs1$13$ ),
    .i1(\picorv32_core/pcpi_rs1$5$ ),
    .sel(\picorv32_core/n555 ),
    .o(\picorv32_core/n558 [9]));  // ../src/picorv32.v(1787)
  binary_mux_s3_w1 \picorv32_core/sel10_b0  (
    .i0(\picorv32_core/mem_rdata_latched [2]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\picorv32_core/n227 [0]),
    .i5(1'b0),
    .i6(\picorv32_core/mem_rdata_latched [2]),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n231 [0]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel10_b1  (
    .i0(\picorv32_core/mem_rdata_latched [3]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\picorv32_core/n227 [1]),
    .i5(1'b0),
    .i6(\picorv32_core/mem_rdata_latched [3]),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n231 [1]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel10_b2  (
    .i0(\picorv32_core/mem_rdata_latched [4]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\picorv32_core/n227 [2]),
    .i5(1'b0),
    .i6(\picorv32_core/mem_rdata_latched [4]),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n231 [2]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel10_b3  (
    .i0(\picorv32_core/mem_rdata_latched [5]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\picorv32_core/n227 [3]),
    .i5(1'b0),
    .i6(\picorv32_core/mem_rdata_latched [5]),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n231 [3]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel10_b4  (
    .i0(\picorv32_core/mem_rdata_latched [6]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\picorv32_core/n227 [4]),
    .i5(1'b0),
    .i6(\picorv32_core/mem_rdata_latched [6]),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n231 [4]));  // ../src/picorv32.v(987)
  and \picorv32_core/sel11_b0/and_b0_1  (\picorv32_core/sel11_b0/B1 , \picorv32_core/mem_rdata_q [7], \picorv32_core/is_sb_sh_sw );
  and \picorv32_core/sel11_b0/and_b0_3  (\picorv32_core/sel11_b0/B3 , \picorv32_core/mem_rdata_q [20], \picorv32_core/n356 );
  or \picorv32_core/sel11_b0/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [0], \picorv32_core/sel11_b0/B1 , \picorv32_core/sel11_b0/B3 );
  and \picorv32_core/sel11_b1/and_b0_1  (\picorv32_core/sel11_b1/B1 , \picorv32_core/mem_rdata_q [8], \picorv32_core/is_sb_sh_sw );
  and \picorv32_core/sel11_b1/and_b0_2  (\picorv32_core/sel11_b1/B2 , \picorv32_core/mem_rdata_q [8], \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/sel11_b1/and_b0_3  (\picorv32_core/sel11_b1/B3 , \picorv32_core/mem_rdata_q [21], \picorv32_core/n356 );
  and \picorv32_core/sel11_b1/and_b0_5  (\picorv32_core/sel11_b1/B5 , \picorv32_core/decoded_imm_uj [1], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b1/or_B1_B2  (\picorv32_core/sel11_b1/or_B1_B2_o , \picorv32_core/sel11_b1/B1 , \picorv32_core/sel11_b1/B2 );
  or \picorv32_core/sel11_b1/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b1/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b1/B3 , \picorv32_core/sel11_b1/B5 );
  or \picorv32_core/sel11_b1/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [1], \picorv32_core/sel11_b1/or_B1_B2_o , \picorv32_core/sel11_b1/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b10/and_b0_1  (\picorv32_core/sel11_b10/B1 , \picorv32_core/mem_rdata_q [30], \picorv32_core/is_sb_sh_sw );
  and \picorv32_core/sel11_b10/and_b0_2  (\picorv32_core/sel11_b10/B2 , \picorv32_core/mem_rdata_q [30], \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/sel11_b10/and_b0_3  (\picorv32_core/sel11_b10/B3 , \picorv32_core/mem_rdata_q [30], \picorv32_core/n356 );
  and \picorv32_core/sel11_b10/and_b0_5  (\picorv32_core/sel11_b10/B5 , \picorv32_core/decoded_imm_uj [10], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b10/or_B1_B2  (\picorv32_core/sel11_b10/or_B1_B2_o , \picorv32_core/sel11_b10/B1 , \picorv32_core/sel11_b10/B2 );
  or \picorv32_core/sel11_b10/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b10/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b10/B3 , \picorv32_core/sel11_b10/B5 );
  or \picorv32_core/sel11_b10/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [10], \picorv32_core/sel11_b10/or_B1_B2_o , \picorv32_core/sel11_b10/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b11/and_b0_1  (\picorv32_core/sel11_b11/B1 , \picorv32_core/mem_rdata_q [31], \picorv32_core/is_sb_sh_sw );
  and \picorv32_core/sel11_b11/and_b0_2  (\picorv32_core/sel11_b11/B2 , \picorv32_core/mem_rdata_q [7], \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/sel11_b11/and_b0_3  (\picorv32_core/sel11_b11/B3 , \picorv32_core/mem_rdata_q [31], \picorv32_core/n356 );
  and \picorv32_core/sel11_b11/and_b0_5  (\picorv32_core/sel11_b11/B5 , \picorv32_core/decoded_imm_uj [11], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b11/or_B1_B2  (\picorv32_core/sel11_b11/or_B1_B2_o , \picorv32_core/sel11_b11/B1 , \picorv32_core/sel11_b11/B2 );
  or \picorv32_core/sel11_b11/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b11/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b11/B5 );
  or \picorv32_core/sel11_b11/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [11], \picorv32_core/sel11_b11/or_B1_B2_o , \picorv32_core/sel11_b11/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b12/and_b0_2  (\picorv32_core/sel11_b12/B2 , \picorv32_core/mem_rdata_q [31], \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/sel11_b12/and_b0_4  (\picorv32_core/sel11_b12/B4 , \picorv32_core/mem_rdata_q [12], \picorv32_core/n473 );
  and \picorv32_core/sel11_b12/and_b0_5  (\picorv32_core/sel11_b12/B5 , \picorv32_core/decoded_imm_uj [12], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b12/or_B1_B2  (\picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b11/B1 , \picorv32_core/sel11_b12/B2 );
  or \picorv32_core/sel11_b12/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b12/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b12/or_B4_B5_o );
  or \picorv32_core/sel11_b12/or_B4_B5  (\picorv32_core/sel11_b12/or_B4_B5_o , \picorv32_core/sel11_b12/B4 , \picorv32_core/sel11_b12/B5 );
  or \picorv32_core/sel11_b12/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [12], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b12/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b13/and_b0_4  (\picorv32_core/sel11_b13/B4 , \picorv32_core/mem_rdata_q [13], \picorv32_core/n473 );
  and \picorv32_core/sel11_b13/and_b0_5  (\picorv32_core/sel11_b13/B5 , \picorv32_core/decoded_imm_uj [13], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b13/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b13/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b13/or_B4_B5_o );
  or \picorv32_core/sel11_b13/or_B4_B5  (\picorv32_core/sel11_b13/or_B4_B5_o , \picorv32_core/sel11_b13/B4 , \picorv32_core/sel11_b13/B5 );
  or \picorv32_core/sel11_b13/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [13], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b13/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b14/and_b0_4  (\picorv32_core/sel11_b14/B4 , \picorv32_core/mem_rdata_q [14], \picorv32_core/n473 );
  and \picorv32_core/sel11_b14/and_b0_5  (\picorv32_core/sel11_b14/B5 , \picorv32_core/decoded_imm_uj [14], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b14/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b14/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b14/or_B4_B5_o );
  or \picorv32_core/sel11_b14/or_B4_B5  (\picorv32_core/sel11_b14/or_B4_B5_o , \picorv32_core/sel11_b14/B4 , \picorv32_core/sel11_b14/B5 );
  or \picorv32_core/sel11_b14/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [14], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b14/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b15/and_b0_4  (\picorv32_core/sel11_b15/B4 , \picorv32_core/mem_rdata_q [15], \picorv32_core/n473 );
  and \picorv32_core/sel11_b15/and_b0_5  (\picorv32_core/sel11_b15/B5 , \picorv32_core/decoded_imm_uj [15], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b15/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b15/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b15/or_B4_B5_o );
  or \picorv32_core/sel11_b15/or_B4_B5  (\picorv32_core/sel11_b15/or_B4_B5_o , \picorv32_core/sel11_b15/B4 , \picorv32_core/sel11_b15/B5 );
  or \picorv32_core/sel11_b15/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [15], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b15/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b16/and_b0_4  (\picorv32_core/sel11_b16/B4 , \picorv32_core/mem_rdata_q [16], \picorv32_core/n473 );
  and \picorv32_core/sel11_b16/and_b0_5  (\picorv32_core/sel11_b16/B5 , \picorv32_core/decoded_imm_uj [16], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b16/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b16/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b16/or_B4_B5_o );
  or \picorv32_core/sel11_b16/or_B4_B5  (\picorv32_core/sel11_b16/or_B4_B5_o , \picorv32_core/sel11_b16/B4 , \picorv32_core/sel11_b16/B5 );
  or \picorv32_core/sel11_b16/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [16], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b16/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b17/and_b0_4  (\picorv32_core/sel11_b17/B4 , \picorv32_core/mem_rdata_q [17], \picorv32_core/n473 );
  and \picorv32_core/sel11_b17/and_b0_5  (\picorv32_core/sel11_b17/B5 , \picorv32_core/decoded_imm_uj [17], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b17/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b17/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b17/or_B4_B5_o );
  or \picorv32_core/sel11_b17/or_B4_B5  (\picorv32_core/sel11_b17/or_B4_B5_o , \picorv32_core/sel11_b17/B4 , \picorv32_core/sel11_b17/B5 );
  or \picorv32_core/sel11_b17/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [17], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b17/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b18/and_b0_4  (\picorv32_core/sel11_b18/B4 , \picorv32_core/mem_rdata_q [18], \picorv32_core/n473 );
  and \picorv32_core/sel11_b18/and_b0_5  (\picorv32_core/sel11_b18/B5 , \picorv32_core/decoded_imm_uj [18], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b18/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b18/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b18/or_B4_B5_o );
  or \picorv32_core/sel11_b18/or_B4_B5  (\picorv32_core/sel11_b18/or_B4_B5_o , \picorv32_core/sel11_b18/B4 , \picorv32_core/sel11_b18/B5 );
  or \picorv32_core/sel11_b18/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [18], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b18/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b19/and_b0_4  (\picorv32_core/sel11_b19/B4 , \picorv32_core/mem_rdata_q [19], \picorv32_core/n473 );
  and \picorv32_core/sel11_b19/and_b0_5  (\picorv32_core/sel11_b19/B5 , \picorv32_core/decoded_imm_uj [19], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b19/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b19/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b19/or_B4_B5_o );
  or \picorv32_core/sel11_b19/or_B4_B5  (\picorv32_core/sel11_b19/or_B4_B5_o , \picorv32_core/sel11_b19/B4 , \picorv32_core/sel11_b19/B5 );
  or \picorv32_core/sel11_b19/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [19], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b19/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b2/and_b0_1  (\picorv32_core/sel11_b2/B1 , \picorv32_core/mem_rdata_q [9], \picorv32_core/is_sb_sh_sw );
  and \picorv32_core/sel11_b2/and_b0_2  (\picorv32_core/sel11_b2/B2 , \picorv32_core/mem_rdata_q [9], \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/sel11_b2/and_b0_3  (\picorv32_core/sel11_b2/B3 , \picorv32_core/mem_rdata_q [22], \picorv32_core/n356 );
  and \picorv32_core/sel11_b2/and_b0_5  (\picorv32_core/sel11_b2/B5 , \picorv32_core/decoded_imm_uj [2], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b2/or_B1_B2  (\picorv32_core/sel11_b2/or_B1_B2_o , \picorv32_core/sel11_b2/B1 , \picorv32_core/sel11_b2/B2 );
  or \picorv32_core/sel11_b2/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b2/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b2/B3 , \picorv32_core/sel11_b2/B5 );
  or \picorv32_core/sel11_b2/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [2], \picorv32_core/sel11_b2/or_B1_B2_o , \picorv32_core/sel11_b2/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b20/and_b0_4  (\picorv32_core/sel11_b20/B4 , \picorv32_core/mem_rdata_q [20], \picorv32_core/n473 );
  and \picorv32_core/sel11_b20/and_b0_5  (\picorv32_core/sel11_b20/B5 , \picorv32_core/decoded_imm_uj [20], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b20/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b20/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b20/or_B4_B5_o );
  or \picorv32_core/sel11_b20/or_B4_B5  (\picorv32_core/sel11_b20/or_B4_B5_o , \picorv32_core/sel11_b20/B4 , \picorv32_core/sel11_b20/B5 );
  or \picorv32_core/sel11_b20/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [20], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b20/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b21/and_b0_4  (\picorv32_core/sel11_b21/B4 , \picorv32_core/mem_rdata_q [21], \picorv32_core/n473 );
  or \picorv32_core/sel11_b21/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b21/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b21/or_B4_B5_o );
  or \picorv32_core/sel11_b21/or_B4_B5  (\picorv32_core/sel11_b21/or_B4_B5_o , \picorv32_core/sel11_b21/B4 , \picorv32_core/sel11_b20/B5 );
  or \picorv32_core/sel11_b21/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [21], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b21/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b22/and_b0_4  (\picorv32_core/sel11_b22/B4 , \picorv32_core/mem_rdata_q [22], \picorv32_core/n473 );
  or \picorv32_core/sel11_b22/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b22/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b22/or_B4_B5_o );
  or \picorv32_core/sel11_b22/or_B4_B5  (\picorv32_core/sel11_b22/or_B4_B5_o , \picorv32_core/sel11_b22/B4 , \picorv32_core/sel11_b20/B5 );
  or \picorv32_core/sel11_b22/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [22], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b22/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b23/and_b0_4  (\picorv32_core/sel11_b23/B4 , \picorv32_core/mem_rdata_q [23], \picorv32_core/n473 );
  or \picorv32_core/sel11_b23/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b23/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b23/or_B4_B5_o );
  or \picorv32_core/sel11_b23/or_B4_B5  (\picorv32_core/sel11_b23/or_B4_B5_o , \picorv32_core/sel11_b23/B4 , \picorv32_core/sel11_b20/B5 );
  or \picorv32_core/sel11_b23/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [23], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b23/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b24/and_b0_4  (\picorv32_core/sel11_b24/B4 , \picorv32_core/mem_rdata_q [24], \picorv32_core/n473 );
  or \picorv32_core/sel11_b24/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b24/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b24/or_B4_B5_o );
  or \picorv32_core/sel11_b24/or_B4_B5  (\picorv32_core/sel11_b24/or_B4_B5_o , \picorv32_core/sel11_b24/B4 , \picorv32_core/sel11_b20/B5 );
  or \picorv32_core/sel11_b24/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [24], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b24/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b25/and_b0_4  (\picorv32_core/sel11_b25/B4 , \picorv32_core/mem_rdata_q [25], \picorv32_core/n473 );
  or \picorv32_core/sel11_b25/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b25/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b25/or_B4_B5_o );
  or \picorv32_core/sel11_b25/or_B4_B5  (\picorv32_core/sel11_b25/or_B4_B5_o , \picorv32_core/sel11_b25/B4 , \picorv32_core/sel11_b20/B5 );
  or \picorv32_core/sel11_b25/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [25], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b25/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b26/and_b0_4  (\picorv32_core/sel11_b26/B4 , \picorv32_core/mem_rdata_q [26], \picorv32_core/n473 );
  or \picorv32_core/sel11_b26/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b26/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b26/or_B4_B5_o );
  or \picorv32_core/sel11_b26/or_B4_B5  (\picorv32_core/sel11_b26/or_B4_B5_o , \picorv32_core/sel11_b26/B4 , \picorv32_core/sel11_b20/B5 );
  or \picorv32_core/sel11_b26/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [26], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b26/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b27/and_b0_4  (\picorv32_core/sel11_b27/B4 , \picorv32_core/mem_rdata_q [27], \picorv32_core/n473 );
  or \picorv32_core/sel11_b27/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b27/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b27/or_B4_B5_o );
  or \picorv32_core/sel11_b27/or_B4_B5  (\picorv32_core/sel11_b27/or_B4_B5_o , \picorv32_core/sel11_b27/B4 , \picorv32_core/sel11_b20/B5 );
  or \picorv32_core/sel11_b27/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [27], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b27/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b28/and_b0_4  (\picorv32_core/sel11_b28/B4 , \picorv32_core/mem_rdata_q [28], \picorv32_core/n473 );
  or \picorv32_core/sel11_b28/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b28/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b28/or_B4_B5_o );
  or \picorv32_core/sel11_b28/or_B4_B5  (\picorv32_core/sel11_b28/or_B4_B5_o , \picorv32_core/sel11_b28/B4 , \picorv32_core/sel11_b20/B5 );
  or \picorv32_core/sel11_b28/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [28], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b28/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b29/and_b0_4  (\picorv32_core/sel11_b29/B4 , \picorv32_core/mem_rdata_q [29], \picorv32_core/n473 );
  or \picorv32_core/sel11_b29/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b29/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b29/or_B4_B5_o );
  or \picorv32_core/sel11_b29/or_B4_B5  (\picorv32_core/sel11_b29/or_B4_B5_o , \picorv32_core/sel11_b29/B4 , \picorv32_core/sel11_b20/B5 );
  or \picorv32_core/sel11_b29/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [29], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b29/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b3/and_b0_1  (\picorv32_core/sel11_b3/B1 , \picorv32_core/mem_rdata_q [10], \picorv32_core/is_sb_sh_sw );
  and \picorv32_core/sel11_b3/and_b0_2  (\picorv32_core/sel11_b3/B2 , \picorv32_core/mem_rdata_q [10], \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/sel11_b3/and_b0_3  (\picorv32_core/sel11_b3/B3 , \picorv32_core/mem_rdata_q [23], \picorv32_core/n356 );
  and \picorv32_core/sel11_b3/and_b0_5  (\picorv32_core/sel11_b3/B5 , \picorv32_core/decoded_imm_uj [3], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b3/or_B1_B2  (\picorv32_core/sel11_b3/or_B1_B2_o , \picorv32_core/sel11_b3/B1 , \picorv32_core/sel11_b3/B2 );
  or \picorv32_core/sel11_b3/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b3/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b3/B3 , \picorv32_core/sel11_b3/B5 );
  or \picorv32_core/sel11_b3/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [3], \picorv32_core/sel11_b3/or_B1_B2_o , \picorv32_core/sel11_b3/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b30/and_b0_4  (\picorv32_core/sel11_b30/B4 , \picorv32_core/mem_rdata_q [30], \picorv32_core/n473 );
  or \picorv32_core/sel11_b30/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b30/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b30/or_B4_B5_o );
  or \picorv32_core/sel11_b30/or_B4_B5  (\picorv32_core/sel11_b30/or_B4_B5_o , \picorv32_core/sel11_b30/B4 , \picorv32_core/sel11_b20/B5 );
  or \picorv32_core/sel11_b30/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [30], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b30/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b31/and_b0_4  (\picorv32_core/sel11_b31/B4 , \picorv32_core/mem_rdata_q [31], \picorv32_core/n473 );
  or \picorv32_core/sel11_b31/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b31/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b11/B3 , \picorv32_core/sel11_b31/or_B4_B5_o );
  or \picorv32_core/sel11_b31/or_B4_B5  (\picorv32_core/sel11_b31/or_B4_B5_o , \picorv32_core/sel11_b31/B4 , \picorv32_core/sel11_b20/B5 );
  or \picorv32_core/sel11_b31/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [31], \picorv32_core/sel11_b12/or_B1_B2_o , \picorv32_core/sel11_b31/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b4/and_b0_1  (\picorv32_core/sel11_b4/B1 , \picorv32_core/mem_rdata_q [11], \picorv32_core/is_sb_sh_sw );
  and \picorv32_core/sel11_b4/and_b0_2  (\picorv32_core/sel11_b4/B2 , \picorv32_core/mem_rdata_q [11], \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/sel11_b4/and_b0_3  (\picorv32_core/sel11_b4/B3 , \picorv32_core/mem_rdata_q [24], \picorv32_core/n356 );
  and \picorv32_core/sel11_b4/and_b0_5  (\picorv32_core/sel11_b4/B5 , \picorv32_core/decoded_imm_uj [4], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b4/or_B1_B2  (\picorv32_core/sel11_b4/or_B1_B2_o , \picorv32_core/sel11_b4/B1 , \picorv32_core/sel11_b4/B2 );
  or \picorv32_core/sel11_b4/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b4/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b4/B3 , \picorv32_core/sel11_b4/B5 );
  or \picorv32_core/sel11_b4/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [4], \picorv32_core/sel11_b4/or_B1_B2_o , \picorv32_core/sel11_b4/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b5/and_b0_1  (\picorv32_core/sel11_b5/B1 , \picorv32_core/mem_rdata_q [25], \picorv32_core/is_sb_sh_sw );
  and \picorv32_core/sel11_b5/and_b0_2  (\picorv32_core/sel11_b5/B2 , \picorv32_core/mem_rdata_q [25], \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/sel11_b5/and_b0_3  (\picorv32_core/sel11_b5/B3 , \picorv32_core/mem_rdata_q [25], \picorv32_core/n356 );
  and \picorv32_core/sel11_b5/and_b0_5  (\picorv32_core/sel11_b5/B5 , \picorv32_core/decoded_imm_uj [5], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b5/or_B1_B2  (\picorv32_core/sel11_b5/or_B1_B2_o , \picorv32_core/sel11_b5/B1 , \picorv32_core/sel11_b5/B2 );
  or \picorv32_core/sel11_b5/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b5/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b5/B3 , \picorv32_core/sel11_b5/B5 );
  or \picorv32_core/sel11_b5/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [5], \picorv32_core/sel11_b5/or_B1_B2_o , \picorv32_core/sel11_b5/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b6/and_b0_1  (\picorv32_core/sel11_b6/B1 , \picorv32_core/mem_rdata_q [26], \picorv32_core/is_sb_sh_sw );
  and \picorv32_core/sel11_b6/and_b0_2  (\picorv32_core/sel11_b6/B2 , \picorv32_core/mem_rdata_q [26], \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/sel11_b6/and_b0_3  (\picorv32_core/sel11_b6/B3 , \picorv32_core/mem_rdata_q [26], \picorv32_core/n356 );
  and \picorv32_core/sel11_b6/and_b0_5  (\picorv32_core/sel11_b6/B5 , \picorv32_core/decoded_imm_uj [6], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b6/or_B1_B2  (\picorv32_core/sel11_b6/or_B1_B2_o , \picorv32_core/sel11_b6/B1 , \picorv32_core/sel11_b6/B2 );
  or \picorv32_core/sel11_b6/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b6/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b6/B3 , \picorv32_core/sel11_b6/B5 );
  or \picorv32_core/sel11_b6/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [6], \picorv32_core/sel11_b6/or_B1_B2_o , \picorv32_core/sel11_b6/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b7/and_b0_1  (\picorv32_core/sel11_b7/B1 , \picorv32_core/mem_rdata_q [27], \picorv32_core/is_sb_sh_sw );
  and \picorv32_core/sel11_b7/and_b0_2  (\picorv32_core/sel11_b7/B2 , \picorv32_core/mem_rdata_q [27], \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/sel11_b7/and_b0_3  (\picorv32_core/sel11_b7/B3 , \picorv32_core/mem_rdata_q [27], \picorv32_core/n356 );
  and \picorv32_core/sel11_b7/and_b0_5  (\picorv32_core/sel11_b7/B5 , \picorv32_core/decoded_imm_uj [7], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b7/or_B1_B2  (\picorv32_core/sel11_b7/or_B1_B2_o , \picorv32_core/sel11_b7/B1 , \picorv32_core/sel11_b7/B2 );
  or \picorv32_core/sel11_b7/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b7/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b7/B3 , \picorv32_core/sel11_b7/B5 );
  or \picorv32_core/sel11_b7/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [7], \picorv32_core/sel11_b7/or_B1_B2_o , \picorv32_core/sel11_b7/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b8/and_b0_1  (\picorv32_core/sel11_b8/B1 , \picorv32_core/mem_rdata_q [28], \picorv32_core/is_sb_sh_sw );
  and \picorv32_core/sel11_b8/and_b0_2  (\picorv32_core/sel11_b8/B2 , \picorv32_core/mem_rdata_q [28], \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/sel11_b8/and_b0_3  (\picorv32_core/sel11_b8/B3 , \picorv32_core/mem_rdata_q [28], \picorv32_core/n356 );
  and \picorv32_core/sel11_b8/and_b0_5  (\picorv32_core/sel11_b8/B5 , \picorv32_core/decoded_imm_uj [8], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b8/or_B1_B2  (\picorv32_core/sel11_b8/or_B1_B2_o , \picorv32_core/sel11_b8/B1 , \picorv32_core/sel11_b8/B2 );
  or \picorv32_core/sel11_b8/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b8/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b8/B3 , \picorv32_core/sel11_b8/B5 );
  or \picorv32_core/sel11_b8/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [8], \picorv32_core/sel11_b8/or_B1_B2_o , \picorv32_core/sel11_b8/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel11_b9/and_b0_1  (\picorv32_core/sel11_b9/B1 , \picorv32_core/mem_rdata_q [29], \picorv32_core/is_sb_sh_sw );
  and \picorv32_core/sel11_b9/and_b0_2  (\picorv32_core/sel11_b9/B2 , \picorv32_core/mem_rdata_q [29], \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/sel11_b9/and_b0_3  (\picorv32_core/sel11_b9/B3 , \picorv32_core/mem_rdata_q [29], \picorv32_core/n356 );
  and \picorv32_core/sel11_b9/and_b0_5  (\picorv32_core/sel11_b9/B5 , \picorv32_core/decoded_imm_uj [9], \picorv32_core/instr_jal );
  or \picorv32_core/sel11_b9/or_B1_B2  (\picorv32_core/sel11_b9/or_B1_B2_o , \picorv32_core/sel11_b9/B1 , \picorv32_core/sel11_b9/B2 );
  or \picorv32_core/sel11_b9/or_B3_or_B4_B5_o  (\picorv32_core/sel11_b9/or_B3_or_B4_B5_o_o , \picorv32_core/sel11_b9/B3 , \picorv32_core/sel11_b9/B5 );
  or \picorv32_core/sel11_b9/or_or_B0_or_B1_B2_o_  (\picorv32_core/n358 [9], \picorv32_core/sel11_b9/or_B1_B2_o , \picorv32_core/sel11_b9/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel12/and_b0_0  (\picorv32_core/sel12/B0 , \picorv32_core/alu_ltu , \picorv32_core/is_sltiu_bltu_sltu );
  and \picorv32_core/sel12/and_b0_1  (\picorv32_core/sel12/B1 , \picorv32_core/alu_lts , \picorv32_core/is_slti_blt_slt );
  and \picorv32_core/sel12/and_b0_2  (\picorv32_core/sel12/B2 , \picorv32_core/n437 , \picorv32_core/instr_bgeu );
  and \picorv32_core/sel12/and_b0_3  (\picorv32_core/sel12/B3 , \picorv32_core/n436 , \picorv32_core/instr_bge );
  or \picorv32_core/sel12/or_B0_or_B1_B2_o  (\picorv32_core/sel12/or_B0_or_B1_B2_o_o , \picorv32_core/sel12/B0 , \picorv32_core/sel12/or_B1_B2_o );
  or \picorv32_core/sel12/or_B1_B2  (\picorv32_core/sel12/or_B1_B2_o , \picorv32_core/sel12/B1 , \picorv32_core/sel12/B2 );
  or \picorv32_core/sel12/or_B3_or_B4_B5_o  (\picorv32_core/sel12/or_B3_or_B4_B5_o_o , \picorv32_core/sel12/B3 , \picorv32_core/sel12/or_B4_B5_o );
  AL_MUX \picorv32_core/sel12/or_B4_B5  (
    .i0(\picorv32_core/instr_bne ),
    .i1(\picorv32_core/instr_beq ),
    .sel(\picorv32_core/alu_eq ),
    .o(\picorv32_core/sel12/or_B4_B5_o ));
  or \picorv32_core/sel12/or_or_B0_or_B1_B2_o_  (\picorv32_core/alu_out_0 , \picorv32_core/sel12/or_B0_or_B1_B2_o_o , \picorv32_core/sel12/or_B3_or_B4_B5_o_o );
  and \picorv32_core/sel13_b0/and_b0_0  (\picorv32_core/sel13_b0/B0 , \picorv32_core/n443 [0], \picorv32_core/n442 );
  and \picorv32_core/sel13_b0/and_b0_1  (\picorv32_core/sel13_b0/B1 , \picorv32_core/n441 [0], \picorv32_core/n440 );
  and \picorv32_core/sel13_b0/and_b0_2  (\picorv32_core/sel13_b0/B2 , \picorv32_core/n439 [0], \picorv32_core/n438 );
  and \picorv32_core/sel13_b0/and_b0_3  (\picorv32_core/sel13_b0/B3 , \picorv32_core/alu_out_0 , \picorv32_core/is_compare );
  and \picorv32_core/sel13_b0/and_b0_4  (\picorv32_core/sel13_b0/B4 , \picorv32_core/alu_add_sub [0], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b0/or_B0_B1  (\picorv32_core/sel13_b0/or_B0_B1_o , \picorv32_core/sel13_b0/B0 , \picorv32_core/sel13_b0/B1 );
  or \picorv32_core/sel13_b0/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b0/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b0/B2 , \picorv32_core/sel13_b0/or_B3_B4_o );
  or \picorv32_core/sel13_b0/or_B3_B4  (\picorv32_core/sel13_b0/or_B3_B4_o , \picorv32_core/sel13_b0/B3 , \picorv32_core/sel13_b0/B4 );
  or \picorv32_core/sel13_b0/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [0], \picorv32_core/sel13_b0/or_B0_B1_o , \picorv32_core/sel13_b0/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b1/and_b0_0  (\picorv32_core/sel13_b1/B0 , \picorv32_core/n443 [1], \picorv32_core/n442 );
  and \picorv32_core/sel13_b1/and_b0_1  (\picorv32_core/sel13_b1/B1 , \picorv32_core/n441 [1], \picorv32_core/n440 );
  and \picorv32_core/sel13_b1/and_b0_2  (\picorv32_core/sel13_b1/B2 , \picorv32_core/n439 [1], \picorv32_core/n438 );
  and \picorv32_core/sel13_b1/and_b0_4  (\picorv32_core/sel13_b1/B4 , \picorv32_core/alu_add_sub [1], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b1/or_B0_B1  (\picorv32_core/sel13_b1/or_B0_B1_o , \picorv32_core/sel13_b1/B0 , \picorv32_core/sel13_b1/B1 );
  or \picorv32_core/sel13_b1/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b1/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b1/B2 , \picorv32_core/sel13_b1/B4 );
  or \picorv32_core/sel13_b1/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [1], \picorv32_core/sel13_b1/or_B0_B1_o , \picorv32_core/sel13_b1/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b10/and_b0_0  (\picorv32_core/sel13_b10/B0 , \picorv32_core/n443 [10], \picorv32_core/n442 );
  and \picorv32_core/sel13_b10/and_b0_1  (\picorv32_core/sel13_b10/B1 , \picorv32_core/n441 [10], \picorv32_core/n440 );
  and \picorv32_core/sel13_b10/and_b0_2  (\picorv32_core/sel13_b10/B2 , \picorv32_core/n439 [10], \picorv32_core/n438 );
  and \picorv32_core/sel13_b10/and_b0_4  (\picorv32_core/sel13_b10/B4 , \picorv32_core/alu_add_sub [10], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b10/or_B0_B1  (\picorv32_core/sel13_b10/or_B0_B1_o , \picorv32_core/sel13_b10/B0 , \picorv32_core/sel13_b10/B1 );
  or \picorv32_core/sel13_b10/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b10/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b10/B2 , \picorv32_core/sel13_b10/B4 );
  or \picorv32_core/sel13_b10/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [10], \picorv32_core/sel13_b10/or_B0_B1_o , \picorv32_core/sel13_b10/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b11/and_b0_0  (\picorv32_core/sel13_b11/B0 , \picorv32_core/n443 [11], \picorv32_core/n442 );
  and \picorv32_core/sel13_b11/and_b0_1  (\picorv32_core/sel13_b11/B1 , \picorv32_core/n441 [11], \picorv32_core/n440 );
  and \picorv32_core/sel13_b11/and_b0_2  (\picorv32_core/sel13_b11/B2 , \picorv32_core/n439 [11], \picorv32_core/n438 );
  and \picorv32_core/sel13_b11/and_b0_4  (\picorv32_core/sel13_b11/B4 , \picorv32_core/alu_add_sub [11], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b11/or_B0_B1  (\picorv32_core/sel13_b11/or_B0_B1_o , \picorv32_core/sel13_b11/B0 , \picorv32_core/sel13_b11/B1 );
  or \picorv32_core/sel13_b11/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b11/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b11/B2 , \picorv32_core/sel13_b11/B4 );
  or \picorv32_core/sel13_b11/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [11], \picorv32_core/sel13_b11/or_B0_B1_o , \picorv32_core/sel13_b11/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b12/and_b0_0  (\picorv32_core/sel13_b12/B0 , \picorv32_core/n443 [12], \picorv32_core/n442 );
  and \picorv32_core/sel13_b12/and_b0_1  (\picorv32_core/sel13_b12/B1 , \picorv32_core/n441 [12], \picorv32_core/n440 );
  and \picorv32_core/sel13_b12/and_b0_2  (\picorv32_core/sel13_b12/B2 , \picorv32_core/n439 [12], \picorv32_core/n438 );
  and \picorv32_core/sel13_b12/and_b0_4  (\picorv32_core/sel13_b12/B4 , \picorv32_core/alu_add_sub [12], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b12/or_B0_B1  (\picorv32_core/sel13_b12/or_B0_B1_o , \picorv32_core/sel13_b12/B0 , \picorv32_core/sel13_b12/B1 );
  or \picorv32_core/sel13_b12/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b12/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b12/B2 , \picorv32_core/sel13_b12/B4 );
  or \picorv32_core/sel13_b12/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [12], \picorv32_core/sel13_b12/or_B0_B1_o , \picorv32_core/sel13_b12/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b13/and_b0_0  (\picorv32_core/sel13_b13/B0 , \picorv32_core/n443 [13], \picorv32_core/n442 );
  and \picorv32_core/sel13_b13/and_b0_1  (\picorv32_core/sel13_b13/B1 , \picorv32_core/n441 [13], \picorv32_core/n440 );
  and \picorv32_core/sel13_b13/and_b0_2  (\picorv32_core/sel13_b13/B2 , \picorv32_core/n439 [13], \picorv32_core/n438 );
  and \picorv32_core/sel13_b13/and_b0_4  (\picorv32_core/sel13_b13/B4 , \picorv32_core/alu_add_sub [13], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b13/or_B0_B1  (\picorv32_core/sel13_b13/or_B0_B1_o , \picorv32_core/sel13_b13/B0 , \picorv32_core/sel13_b13/B1 );
  or \picorv32_core/sel13_b13/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b13/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b13/B2 , \picorv32_core/sel13_b13/B4 );
  or \picorv32_core/sel13_b13/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [13], \picorv32_core/sel13_b13/or_B0_B1_o , \picorv32_core/sel13_b13/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b14/and_b0_0  (\picorv32_core/sel13_b14/B0 , \picorv32_core/n443 [14], \picorv32_core/n442 );
  and \picorv32_core/sel13_b14/and_b0_1  (\picorv32_core/sel13_b14/B1 , \picorv32_core/n441 [14], \picorv32_core/n440 );
  and \picorv32_core/sel13_b14/and_b0_2  (\picorv32_core/sel13_b14/B2 , \picorv32_core/n439 [14], \picorv32_core/n438 );
  and \picorv32_core/sel13_b14/and_b0_4  (\picorv32_core/sel13_b14/B4 , \picorv32_core/alu_add_sub [14], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b14/or_B0_B1  (\picorv32_core/sel13_b14/or_B0_B1_o , \picorv32_core/sel13_b14/B0 , \picorv32_core/sel13_b14/B1 );
  or \picorv32_core/sel13_b14/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b14/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b14/B2 , \picorv32_core/sel13_b14/B4 );
  or \picorv32_core/sel13_b14/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [14], \picorv32_core/sel13_b14/or_B0_B1_o , \picorv32_core/sel13_b14/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b15/and_b0_0  (\picorv32_core/sel13_b15/B0 , \picorv32_core/n443 [15], \picorv32_core/n442 );
  and \picorv32_core/sel13_b15/and_b0_1  (\picorv32_core/sel13_b15/B1 , \picorv32_core/n441 [15], \picorv32_core/n440 );
  and \picorv32_core/sel13_b15/and_b0_2  (\picorv32_core/sel13_b15/B2 , \picorv32_core/n439 [15], \picorv32_core/n438 );
  and \picorv32_core/sel13_b15/and_b0_4  (\picorv32_core/sel13_b15/B4 , \picorv32_core/alu_add_sub [15], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b15/or_B0_B1  (\picorv32_core/sel13_b15/or_B0_B1_o , \picorv32_core/sel13_b15/B0 , \picorv32_core/sel13_b15/B1 );
  or \picorv32_core/sel13_b15/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b15/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b15/B2 , \picorv32_core/sel13_b15/B4 );
  or \picorv32_core/sel13_b15/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [15], \picorv32_core/sel13_b15/or_B0_B1_o , \picorv32_core/sel13_b15/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b16/and_b0_0  (\picorv32_core/sel13_b16/B0 , \picorv32_core/n443 [16], \picorv32_core/n442 );
  and \picorv32_core/sel13_b16/and_b0_1  (\picorv32_core/sel13_b16/B1 , \picorv32_core/n441 [16], \picorv32_core/n440 );
  and \picorv32_core/sel13_b16/and_b0_2  (\picorv32_core/sel13_b16/B2 , \picorv32_core/n439 [16], \picorv32_core/n438 );
  and \picorv32_core/sel13_b16/and_b0_4  (\picorv32_core/sel13_b16/B4 , \picorv32_core/alu_add_sub [16], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b16/or_B0_B1  (\picorv32_core/sel13_b16/or_B0_B1_o , \picorv32_core/sel13_b16/B0 , \picorv32_core/sel13_b16/B1 );
  or \picorv32_core/sel13_b16/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b16/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b16/B2 , \picorv32_core/sel13_b16/B4 );
  or \picorv32_core/sel13_b16/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [16], \picorv32_core/sel13_b16/or_B0_B1_o , \picorv32_core/sel13_b16/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b17/and_b0_0  (\picorv32_core/sel13_b17/B0 , \picorv32_core/n443 [17], \picorv32_core/n442 );
  and \picorv32_core/sel13_b17/and_b0_1  (\picorv32_core/sel13_b17/B1 , \picorv32_core/n441 [17], \picorv32_core/n440 );
  and \picorv32_core/sel13_b17/and_b0_2  (\picorv32_core/sel13_b17/B2 , \picorv32_core/n439 [17], \picorv32_core/n438 );
  and \picorv32_core/sel13_b17/and_b0_4  (\picorv32_core/sel13_b17/B4 , \picorv32_core/alu_add_sub [17], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b17/or_B0_B1  (\picorv32_core/sel13_b17/or_B0_B1_o , \picorv32_core/sel13_b17/B0 , \picorv32_core/sel13_b17/B1 );
  or \picorv32_core/sel13_b17/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b17/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b17/B2 , \picorv32_core/sel13_b17/B4 );
  or \picorv32_core/sel13_b17/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [17], \picorv32_core/sel13_b17/or_B0_B1_o , \picorv32_core/sel13_b17/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b18/and_b0_0  (\picorv32_core/sel13_b18/B0 , \picorv32_core/n443 [18], \picorv32_core/n442 );
  and \picorv32_core/sel13_b18/and_b0_1  (\picorv32_core/sel13_b18/B1 , \picorv32_core/n441 [18], \picorv32_core/n440 );
  and \picorv32_core/sel13_b18/and_b0_2  (\picorv32_core/sel13_b18/B2 , \picorv32_core/n439 [18], \picorv32_core/n438 );
  and \picorv32_core/sel13_b18/and_b0_4  (\picorv32_core/sel13_b18/B4 , \picorv32_core/alu_add_sub [18], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b18/or_B0_B1  (\picorv32_core/sel13_b18/or_B0_B1_o , \picorv32_core/sel13_b18/B0 , \picorv32_core/sel13_b18/B1 );
  or \picorv32_core/sel13_b18/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b18/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b18/B2 , \picorv32_core/sel13_b18/B4 );
  or \picorv32_core/sel13_b18/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [18], \picorv32_core/sel13_b18/or_B0_B1_o , \picorv32_core/sel13_b18/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b19/and_b0_0  (\picorv32_core/sel13_b19/B0 , \picorv32_core/n443 [19], \picorv32_core/n442 );
  and \picorv32_core/sel13_b19/and_b0_1  (\picorv32_core/sel13_b19/B1 , \picorv32_core/n441 [19], \picorv32_core/n440 );
  and \picorv32_core/sel13_b19/and_b0_2  (\picorv32_core/sel13_b19/B2 , \picorv32_core/n439 [19], \picorv32_core/n438 );
  and \picorv32_core/sel13_b19/and_b0_4  (\picorv32_core/sel13_b19/B4 , \picorv32_core/alu_add_sub [19], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b19/or_B0_B1  (\picorv32_core/sel13_b19/or_B0_B1_o , \picorv32_core/sel13_b19/B0 , \picorv32_core/sel13_b19/B1 );
  or \picorv32_core/sel13_b19/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b19/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b19/B2 , \picorv32_core/sel13_b19/B4 );
  or \picorv32_core/sel13_b19/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [19], \picorv32_core/sel13_b19/or_B0_B1_o , \picorv32_core/sel13_b19/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b2/and_b0_0  (\picorv32_core/sel13_b2/B0 , \picorv32_core/n443 [2], \picorv32_core/n442 );
  and \picorv32_core/sel13_b2/and_b0_1  (\picorv32_core/sel13_b2/B1 , \picorv32_core/n441 [2], \picorv32_core/n440 );
  and \picorv32_core/sel13_b2/and_b0_2  (\picorv32_core/sel13_b2/B2 , \picorv32_core/n439 [2], \picorv32_core/n438 );
  and \picorv32_core/sel13_b2/and_b0_4  (\picorv32_core/sel13_b2/B4 , \picorv32_core/alu_add_sub [2], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b2/or_B0_B1  (\picorv32_core/sel13_b2/or_B0_B1_o , \picorv32_core/sel13_b2/B0 , \picorv32_core/sel13_b2/B1 );
  or \picorv32_core/sel13_b2/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b2/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b2/B2 , \picorv32_core/sel13_b2/B4 );
  or \picorv32_core/sel13_b2/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [2], \picorv32_core/sel13_b2/or_B0_B1_o , \picorv32_core/sel13_b2/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b20/and_b0_0  (\picorv32_core/sel13_b20/B0 , \picorv32_core/n443 [20], \picorv32_core/n442 );
  and \picorv32_core/sel13_b20/and_b0_1  (\picorv32_core/sel13_b20/B1 , \picorv32_core/n441 [20], \picorv32_core/n440 );
  and \picorv32_core/sel13_b20/and_b0_2  (\picorv32_core/sel13_b20/B2 , \picorv32_core/n439 [20], \picorv32_core/n438 );
  and \picorv32_core/sel13_b20/and_b0_4  (\picorv32_core/sel13_b20/B4 , \picorv32_core/alu_add_sub [20], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b20/or_B0_B1  (\picorv32_core/sel13_b20/or_B0_B1_o , \picorv32_core/sel13_b20/B0 , \picorv32_core/sel13_b20/B1 );
  or \picorv32_core/sel13_b20/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b20/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b20/B2 , \picorv32_core/sel13_b20/B4 );
  or \picorv32_core/sel13_b20/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [20], \picorv32_core/sel13_b20/or_B0_B1_o , \picorv32_core/sel13_b20/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b21/and_b0_0  (\picorv32_core/sel13_b21/B0 , \picorv32_core/n443 [21], \picorv32_core/n442 );
  and \picorv32_core/sel13_b21/and_b0_1  (\picorv32_core/sel13_b21/B1 , \picorv32_core/n441 [21], \picorv32_core/n440 );
  and \picorv32_core/sel13_b21/and_b0_2  (\picorv32_core/sel13_b21/B2 , \picorv32_core/n439 [21], \picorv32_core/n438 );
  and \picorv32_core/sel13_b21/and_b0_4  (\picorv32_core/sel13_b21/B4 , \picorv32_core/alu_add_sub [21], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b21/or_B0_B1  (\picorv32_core/sel13_b21/or_B0_B1_o , \picorv32_core/sel13_b21/B0 , \picorv32_core/sel13_b21/B1 );
  or \picorv32_core/sel13_b21/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b21/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b21/B2 , \picorv32_core/sel13_b21/B4 );
  or \picorv32_core/sel13_b21/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [21], \picorv32_core/sel13_b21/or_B0_B1_o , \picorv32_core/sel13_b21/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b22/and_b0_0  (\picorv32_core/sel13_b22/B0 , \picorv32_core/n443 [22], \picorv32_core/n442 );
  and \picorv32_core/sel13_b22/and_b0_1  (\picorv32_core/sel13_b22/B1 , \picorv32_core/n441 [22], \picorv32_core/n440 );
  and \picorv32_core/sel13_b22/and_b0_2  (\picorv32_core/sel13_b22/B2 , \picorv32_core/n439 [22], \picorv32_core/n438 );
  and \picorv32_core/sel13_b22/and_b0_4  (\picorv32_core/sel13_b22/B4 , \picorv32_core/alu_add_sub [22], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b22/or_B0_B1  (\picorv32_core/sel13_b22/or_B0_B1_o , \picorv32_core/sel13_b22/B0 , \picorv32_core/sel13_b22/B1 );
  or \picorv32_core/sel13_b22/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b22/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b22/B2 , \picorv32_core/sel13_b22/B4 );
  or \picorv32_core/sel13_b22/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [22], \picorv32_core/sel13_b22/or_B0_B1_o , \picorv32_core/sel13_b22/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b23/and_b0_0  (\picorv32_core/sel13_b23/B0 , \picorv32_core/n443 [23], \picorv32_core/n442 );
  and \picorv32_core/sel13_b23/and_b0_1  (\picorv32_core/sel13_b23/B1 , \picorv32_core/n441 [23], \picorv32_core/n440 );
  and \picorv32_core/sel13_b23/and_b0_2  (\picorv32_core/sel13_b23/B2 , \picorv32_core/n439 [23], \picorv32_core/n438 );
  and \picorv32_core/sel13_b23/and_b0_4  (\picorv32_core/sel13_b23/B4 , \picorv32_core/alu_add_sub [23], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b23/or_B0_B1  (\picorv32_core/sel13_b23/or_B0_B1_o , \picorv32_core/sel13_b23/B0 , \picorv32_core/sel13_b23/B1 );
  or \picorv32_core/sel13_b23/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b23/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b23/B2 , \picorv32_core/sel13_b23/B4 );
  or \picorv32_core/sel13_b23/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [23], \picorv32_core/sel13_b23/or_B0_B1_o , \picorv32_core/sel13_b23/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b24/and_b0_0  (\picorv32_core/sel13_b24/B0 , \picorv32_core/n443 [24], \picorv32_core/n442 );
  and \picorv32_core/sel13_b24/and_b0_1  (\picorv32_core/sel13_b24/B1 , \picorv32_core/n441 [24], \picorv32_core/n440 );
  and \picorv32_core/sel13_b24/and_b0_2  (\picorv32_core/sel13_b24/B2 , \picorv32_core/n439 [24], \picorv32_core/n438 );
  and \picorv32_core/sel13_b24/and_b0_4  (\picorv32_core/sel13_b24/B4 , \picorv32_core/alu_add_sub [24], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b24/or_B0_B1  (\picorv32_core/sel13_b24/or_B0_B1_o , \picorv32_core/sel13_b24/B0 , \picorv32_core/sel13_b24/B1 );
  or \picorv32_core/sel13_b24/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b24/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b24/B2 , \picorv32_core/sel13_b24/B4 );
  or \picorv32_core/sel13_b24/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [24], \picorv32_core/sel13_b24/or_B0_B1_o , \picorv32_core/sel13_b24/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b25/and_b0_0  (\picorv32_core/sel13_b25/B0 , \picorv32_core/n443 [25], \picorv32_core/n442 );
  and \picorv32_core/sel13_b25/and_b0_1  (\picorv32_core/sel13_b25/B1 , \picorv32_core/n441 [25], \picorv32_core/n440 );
  and \picorv32_core/sel13_b25/and_b0_2  (\picorv32_core/sel13_b25/B2 , \picorv32_core/n439 [25], \picorv32_core/n438 );
  and \picorv32_core/sel13_b25/and_b0_4  (\picorv32_core/sel13_b25/B4 , \picorv32_core/alu_add_sub [25], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b25/or_B0_B1  (\picorv32_core/sel13_b25/or_B0_B1_o , \picorv32_core/sel13_b25/B0 , \picorv32_core/sel13_b25/B1 );
  or \picorv32_core/sel13_b25/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b25/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b25/B2 , \picorv32_core/sel13_b25/B4 );
  or \picorv32_core/sel13_b25/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [25], \picorv32_core/sel13_b25/or_B0_B1_o , \picorv32_core/sel13_b25/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b26/and_b0_0  (\picorv32_core/sel13_b26/B0 , \picorv32_core/n443 [26], \picorv32_core/n442 );
  and \picorv32_core/sel13_b26/and_b0_1  (\picorv32_core/sel13_b26/B1 , \picorv32_core/n441 [26], \picorv32_core/n440 );
  and \picorv32_core/sel13_b26/and_b0_2  (\picorv32_core/sel13_b26/B2 , \picorv32_core/n439 [26], \picorv32_core/n438 );
  and \picorv32_core/sel13_b26/and_b0_4  (\picorv32_core/sel13_b26/B4 , \picorv32_core/alu_add_sub [26], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b26/or_B0_B1  (\picorv32_core/sel13_b26/or_B0_B1_o , \picorv32_core/sel13_b26/B0 , \picorv32_core/sel13_b26/B1 );
  or \picorv32_core/sel13_b26/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b26/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b26/B2 , \picorv32_core/sel13_b26/B4 );
  or \picorv32_core/sel13_b26/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [26], \picorv32_core/sel13_b26/or_B0_B1_o , \picorv32_core/sel13_b26/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b27/and_b0_0  (\picorv32_core/sel13_b27/B0 , \picorv32_core/n443 [27], \picorv32_core/n442 );
  and \picorv32_core/sel13_b27/and_b0_1  (\picorv32_core/sel13_b27/B1 , \picorv32_core/n441 [27], \picorv32_core/n440 );
  and \picorv32_core/sel13_b27/and_b0_2  (\picorv32_core/sel13_b27/B2 , \picorv32_core/n439 [27], \picorv32_core/n438 );
  and \picorv32_core/sel13_b27/and_b0_4  (\picorv32_core/sel13_b27/B4 , \picorv32_core/alu_add_sub [27], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b27/or_B0_B1  (\picorv32_core/sel13_b27/or_B0_B1_o , \picorv32_core/sel13_b27/B0 , \picorv32_core/sel13_b27/B1 );
  or \picorv32_core/sel13_b27/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b27/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b27/B2 , \picorv32_core/sel13_b27/B4 );
  or \picorv32_core/sel13_b27/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [27], \picorv32_core/sel13_b27/or_B0_B1_o , \picorv32_core/sel13_b27/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b28/and_b0_0  (\picorv32_core/sel13_b28/B0 , \picorv32_core/n443 [28], \picorv32_core/n442 );
  and \picorv32_core/sel13_b28/and_b0_1  (\picorv32_core/sel13_b28/B1 , \picorv32_core/n441 [28], \picorv32_core/n440 );
  and \picorv32_core/sel13_b28/and_b0_2  (\picorv32_core/sel13_b28/B2 , \picorv32_core/n439 [28], \picorv32_core/n438 );
  and \picorv32_core/sel13_b28/and_b0_4  (\picorv32_core/sel13_b28/B4 , \picorv32_core/alu_add_sub [28], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b28/or_B0_B1  (\picorv32_core/sel13_b28/or_B0_B1_o , \picorv32_core/sel13_b28/B0 , \picorv32_core/sel13_b28/B1 );
  or \picorv32_core/sel13_b28/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b28/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b28/B2 , \picorv32_core/sel13_b28/B4 );
  or \picorv32_core/sel13_b28/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [28], \picorv32_core/sel13_b28/or_B0_B1_o , \picorv32_core/sel13_b28/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b29/and_b0_0  (\picorv32_core/sel13_b29/B0 , \picorv32_core/n443 [29], \picorv32_core/n442 );
  and \picorv32_core/sel13_b29/and_b0_1  (\picorv32_core/sel13_b29/B1 , \picorv32_core/n441 [29], \picorv32_core/n440 );
  and \picorv32_core/sel13_b29/and_b0_2  (\picorv32_core/sel13_b29/B2 , \picorv32_core/n439 [29], \picorv32_core/n438 );
  and \picorv32_core/sel13_b29/and_b0_4  (\picorv32_core/sel13_b29/B4 , \picorv32_core/alu_add_sub [29], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b29/or_B0_B1  (\picorv32_core/sel13_b29/or_B0_B1_o , \picorv32_core/sel13_b29/B0 , \picorv32_core/sel13_b29/B1 );
  or \picorv32_core/sel13_b29/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b29/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b29/B2 , \picorv32_core/sel13_b29/B4 );
  or \picorv32_core/sel13_b29/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [29], \picorv32_core/sel13_b29/or_B0_B1_o , \picorv32_core/sel13_b29/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b3/and_b0_0  (\picorv32_core/sel13_b3/B0 , \picorv32_core/n443 [3], \picorv32_core/n442 );
  and \picorv32_core/sel13_b3/and_b0_1  (\picorv32_core/sel13_b3/B1 , \picorv32_core/n441 [3], \picorv32_core/n440 );
  and \picorv32_core/sel13_b3/and_b0_2  (\picorv32_core/sel13_b3/B2 , \picorv32_core/n439 [3], \picorv32_core/n438 );
  and \picorv32_core/sel13_b3/and_b0_4  (\picorv32_core/sel13_b3/B4 , \picorv32_core/alu_add_sub [3], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b3/or_B0_B1  (\picorv32_core/sel13_b3/or_B0_B1_o , \picorv32_core/sel13_b3/B0 , \picorv32_core/sel13_b3/B1 );
  or \picorv32_core/sel13_b3/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b3/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b3/B2 , \picorv32_core/sel13_b3/B4 );
  or \picorv32_core/sel13_b3/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [3], \picorv32_core/sel13_b3/or_B0_B1_o , \picorv32_core/sel13_b3/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b30/and_b0_0  (\picorv32_core/sel13_b30/B0 , \picorv32_core/n443 [30], \picorv32_core/n442 );
  and \picorv32_core/sel13_b30/and_b0_1  (\picorv32_core/sel13_b30/B1 , \picorv32_core/n441 [30], \picorv32_core/n440 );
  and \picorv32_core/sel13_b30/and_b0_2  (\picorv32_core/sel13_b30/B2 , \picorv32_core/n439 [30], \picorv32_core/n438 );
  and \picorv32_core/sel13_b30/and_b0_4  (\picorv32_core/sel13_b30/B4 , \picorv32_core/alu_add_sub [30], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b30/or_B0_B1  (\picorv32_core/sel13_b30/or_B0_B1_o , \picorv32_core/sel13_b30/B0 , \picorv32_core/sel13_b30/B1 );
  or \picorv32_core/sel13_b30/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b30/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b30/B2 , \picorv32_core/sel13_b30/B4 );
  or \picorv32_core/sel13_b30/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [30], \picorv32_core/sel13_b30/or_B0_B1_o , \picorv32_core/sel13_b30/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b31/and_b0_0  (\picorv32_core/sel13_b31/B0 , \picorv32_core/n443 [31], \picorv32_core/n442 );
  and \picorv32_core/sel13_b31/and_b0_1  (\picorv32_core/sel13_b31/B1 , \picorv32_core/n441 [31], \picorv32_core/n440 );
  and \picorv32_core/sel13_b31/and_b0_2  (\picorv32_core/sel13_b31/B2 , \picorv32_core/n439 [31], \picorv32_core/n438 );
  and \picorv32_core/sel13_b31/and_b0_4  (\picorv32_core/sel13_b31/B4 , \picorv32_core/alu_add_sub [31], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b31/or_B0_B1  (\picorv32_core/sel13_b31/or_B0_B1_o , \picorv32_core/sel13_b31/B0 , \picorv32_core/sel13_b31/B1 );
  or \picorv32_core/sel13_b31/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b31/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b31/B2 , \picorv32_core/sel13_b31/B4 );
  or \picorv32_core/sel13_b31/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [31], \picorv32_core/sel13_b31/or_B0_B1_o , \picorv32_core/sel13_b31/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b4/and_b0_0  (\picorv32_core/sel13_b4/B0 , \picorv32_core/n443 [4], \picorv32_core/n442 );
  and \picorv32_core/sel13_b4/and_b0_1  (\picorv32_core/sel13_b4/B1 , \picorv32_core/n441 [4], \picorv32_core/n440 );
  and \picorv32_core/sel13_b4/and_b0_2  (\picorv32_core/sel13_b4/B2 , \picorv32_core/n439 [4], \picorv32_core/n438 );
  and \picorv32_core/sel13_b4/and_b0_4  (\picorv32_core/sel13_b4/B4 , \picorv32_core/alu_add_sub [4], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b4/or_B0_B1  (\picorv32_core/sel13_b4/or_B0_B1_o , \picorv32_core/sel13_b4/B0 , \picorv32_core/sel13_b4/B1 );
  or \picorv32_core/sel13_b4/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b4/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b4/B2 , \picorv32_core/sel13_b4/B4 );
  or \picorv32_core/sel13_b4/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [4], \picorv32_core/sel13_b4/or_B0_B1_o , \picorv32_core/sel13_b4/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b5/and_b0_0  (\picorv32_core/sel13_b5/B0 , \picorv32_core/n443 [5], \picorv32_core/n442 );
  and \picorv32_core/sel13_b5/and_b0_1  (\picorv32_core/sel13_b5/B1 , \picorv32_core/n441 [5], \picorv32_core/n440 );
  and \picorv32_core/sel13_b5/and_b0_2  (\picorv32_core/sel13_b5/B2 , \picorv32_core/n439 [5], \picorv32_core/n438 );
  and \picorv32_core/sel13_b5/and_b0_4  (\picorv32_core/sel13_b5/B4 , \picorv32_core/alu_add_sub [5], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b5/or_B0_B1  (\picorv32_core/sel13_b5/or_B0_B1_o , \picorv32_core/sel13_b5/B0 , \picorv32_core/sel13_b5/B1 );
  or \picorv32_core/sel13_b5/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b5/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b5/B2 , \picorv32_core/sel13_b5/B4 );
  or \picorv32_core/sel13_b5/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [5], \picorv32_core/sel13_b5/or_B0_B1_o , \picorv32_core/sel13_b5/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b6/and_b0_0  (\picorv32_core/sel13_b6/B0 , \picorv32_core/n443 [6], \picorv32_core/n442 );
  and \picorv32_core/sel13_b6/and_b0_1  (\picorv32_core/sel13_b6/B1 , \picorv32_core/n441 [6], \picorv32_core/n440 );
  and \picorv32_core/sel13_b6/and_b0_2  (\picorv32_core/sel13_b6/B2 , \picorv32_core/n439 [6], \picorv32_core/n438 );
  and \picorv32_core/sel13_b6/and_b0_4  (\picorv32_core/sel13_b6/B4 , \picorv32_core/alu_add_sub [6], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b6/or_B0_B1  (\picorv32_core/sel13_b6/or_B0_B1_o , \picorv32_core/sel13_b6/B0 , \picorv32_core/sel13_b6/B1 );
  or \picorv32_core/sel13_b6/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b6/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b6/B2 , \picorv32_core/sel13_b6/B4 );
  or \picorv32_core/sel13_b6/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [6], \picorv32_core/sel13_b6/or_B0_B1_o , \picorv32_core/sel13_b6/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b7/and_b0_0  (\picorv32_core/sel13_b7/B0 , \picorv32_core/n443 [7], \picorv32_core/n442 );
  and \picorv32_core/sel13_b7/and_b0_1  (\picorv32_core/sel13_b7/B1 , \picorv32_core/n441 [7], \picorv32_core/n440 );
  and \picorv32_core/sel13_b7/and_b0_2  (\picorv32_core/sel13_b7/B2 , \picorv32_core/n439 [7], \picorv32_core/n438 );
  and \picorv32_core/sel13_b7/and_b0_4  (\picorv32_core/sel13_b7/B4 , \picorv32_core/alu_add_sub [7], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b7/or_B0_B1  (\picorv32_core/sel13_b7/or_B0_B1_o , \picorv32_core/sel13_b7/B0 , \picorv32_core/sel13_b7/B1 );
  or \picorv32_core/sel13_b7/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b7/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b7/B2 , \picorv32_core/sel13_b7/B4 );
  or \picorv32_core/sel13_b7/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [7], \picorv32_core/sel13_b7/or_B0_B1_o , \picorv32_core/sel13_b7/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b8/and_b0_0  (\picorv32_core/sel13_b8/B0 , \picorv32_core/n443 [8], \picorv32_core/n442 );
  and \picorv32_core/sel13_b8/and_b0_1  (\picorv32_core/sel13_b8/B1 , \picorv32_core/n441 [8], \picorv32_core/n440 );
  and \picorv32_core/sel13_b8/and_b0_2  (\picorv32_core/sel13_b8/B2 , \picorv32_core/n439 [8], \picorv32_core/n438 );
  and \picorv32_core/sel13_b8/and_b0_4  (\picorv32_core/sel13_b8/B4 , \picorv32_core/alu_add_sub [8], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b8/or_B0_B1  (\picorv32_core/sel13_b8/or_B0_B1_o , \picorv32_core/sel13_b8/B0 , \picorv32_core/sel13_b8/B1 );
  or \picorv32_core/sel13_b8/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b8/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b8/B2 , \picorv32_core/sel13_b8/B4 );
  or \picorv32_core/sel13_b8/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [8], \picorv32_core/sel13_b8/or_B0_B1_o , \picorv32_core/sel13_b8/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel13_b9/and_b0_0  (\picorv32_core/sel13_b9/B0 , \picorv32_core/n443 [9], \picorv32_core/n442 );
  and \picorv32_core/sel13_b9/and_b0_1  (\picorv32_core/sel13_b9/B1 , \picorv32_core/n441 [9], \picorv32_core/n440 );
  and \picorv32_core/sel13_b9/and_b0_2  (\picorv32_core/sel13_b9/B2 , \picorv32_core/n439 [9], \picorv32_core/n438 );
  and \picorv32_core/sel13_b9/and_b0_4  (\picorv32_core/sel13_b9/B4 , \picorv32_core/alu_add_sub [9], \picorv32_core/is_lui_auipc_jal_jalr_addi_add_sub );
  or \picorv32_core/sel13_b9/or_B0_B1  (\picorv32_core/sel13_b9/or_B0_B1_o , \picorv32_core/sel13_b9/B0 , \picorv32_core/sel13_b9/B1 );
  or \picorv32_core/sel13_b9/or_B2_or_B3_B4_o  (\picorv32_core/sel13_b9/or_B2_or_B3_B4_o_o , \picorv32_core/sel13_b9/B2 , \picorv32_core/sel13_b9/B4 );
  or \picorv32_core/sel13_b9/or_or_B0_B1_o_or_B2_  (\picorv32_core/alu_out [9], \picorv32_core/sel13_b9/or_B0_B1_o , \picorv32_core/sel13_b9/or_B2_or_B3_B4_o_o );
  AL_MUX \picorv32_core/sel14_b0  (
    .i0(\picorv32_core/n453 [0]),
    .i1(\picorv32_core/n450 [0]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [0]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b1  (
    .i0(\picorv32_core/n453 [1]),
    .i1(\picorv32_core/n450 [1]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [1]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b10  (
    .i0(\picorv32_core/n453 [10]),
    .i1(\picorv32_core/n450 [10]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [10]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b11  (
    .i0(\picorv32_core/n453 [11]),
    .i1(\picorv32_core/n450 [11]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [11]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b12  (
    .i0(\picorv32_core/n453 [12]),
    .i1(\picorv32_core/n450 [12]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [12]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b13  (
    .i0(\picorv32_core/n453 [13]),
    .i1(\picorv32_core/n450 [13]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [13]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b14  (
    .i0(\picorv32_core/n453 [14]),
    .i1(\picorv32_core/n450 [14]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [14]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b15  (
    .i0(\picorv32_core/n453 [15]),
    .i1(\picorv32_core/n450 [15]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [15]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b16  (
    .i0(\picorv32_core/n453 [16]),
    .i1(\picorv32_core/n450 [16]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [16]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b17  (
    .i0(\picorv32_core/n453 [17]),
    .i1(\picorv32_core/n450 [17]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [17]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b18  (
    .i0(\picorv32_core/n453 [18]),
    .i1(\picorv32_core/n450 [18]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [18]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b19  (
    .i0(\picorv32_core/n453 [19]),
    .i1(\picorv32_core/n450 [19]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [19]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b2  (
    .i0(\picorv32_core/n453 [2]),
    .i1(\picorv32_core/n450 [2]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [2]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b20  (
    .i0(\picorv32_core/n453 [20]),
    .i1(\picorv32_core/n450 [20]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [20]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b21  (
    .i0(\picorv32_core/n453 [21]),
    .i1(\picorv32_core/n450 [21]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [21]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b22  (
    .i0(\picorv32_core/n453 [22]),
    .i1(\picorv32_core/n450 [22]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [22]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b23  (
    .i0(\picorv32_core/n453 [23]),
    .i1(\picorv32_core/n450 [23]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [23]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b24  (
    .i0(\picorv32_core/n453 [24]),
    .i1(\picorv32_core/n450 [24]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [24]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b25  (
    .i0(\picorv32_core/n453 [25]),
    .i1(\picorv32_core/n450 [25]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [25]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b26  (
    .i0(\picorv32_core/n453 [26]),
    .i1(\picorv32_core/n450 [26]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [26]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b27  (
    .i0(\picorv32_core/n453 [27]),
    .i1(\picorv32_core/n450 [27]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [27]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b28  (
    .i0(\picorv32_core/n453 [28]),
    .i1(\picorv32_core/n450 [28]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [28]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b29  (
    .i0(\picorv32_core/n453 [29]),
    .i1(\picorv32_core/n450 [29]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [29]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b3  (
    .i0(\picorv32_core/n453 [3]),
    .i1(\picorv32_core/n450 [3]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [3]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b30  (
    .i0(\picorv32_core/n453 [30]),
    .i1(\picorv32_core/n450 [30]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [30]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b31  (
    .i0(\picorv32_core/n453 [31]),
    .i1(\picorv32_core/n450 [31]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [31]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b4  (
    .i0(\picorv32_core/n453 [4]),
    .i1(\picorv32_core/n450 [4]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [4]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b5  (
    .i0(\picorv32_core/n453 [5]),
    .i1(\picorv32_core/n450 [5]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [5]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b6  (
    .i0(\picorv32_core/n453 [6]),
    .i1(\picorv32_core/n450 [6]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [6]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b7  (
    .i0(\picorv32_core/n453 [7]),
    .i1(\picorv32_core/n450 [7]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [7]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b8  (
    .i0(\picorv32_core/n453 [8]),
    .i1(\picorv32_core/n450 [8]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [8]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel14_b9  (
    .i0(\picorv32_core/n453 [9]),
    .i1(\picorv32_core/n450 [9]),
    .sel(\picorv32_core/latched_branch ),
    .o(\picorv32_core/n455 [9]));  // ../src/picorv32.v(1285)
  AL_MUX \picorv32_core/sel15_b0  (
    .i0(\picorv32_core/reg_next_pc [0]),
    .i1(\picorv32_core/n453 [0]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [0]));
  and \picorv32_core/sel15_b0_sel_is_3  (\picorv32_core/sel15_b0_sel_is_3_o , \picorv32_core/latched_branch , \picorv32_core/latched_store );
  AL_MUX \picorv32_core/sel15_b1  (
    .i0(\picorv32_core/reg_next_pc [1]),
    .i1(\picorv32_core/n453 [1]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [1]));
  AL_MUX \picorv32_core/sel15_b10  (
    .i0(\picorv32_core/reg_next_pc [10]),
    .i1(\picorv32_core/n453 [10]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [10]));
  AL_MUX \picorv32_core/sel15_b11  (
    .i0(\picorv32_core/reg_next_pc [11]),
    .i1(\picorv32_core/n453 [11]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [11]));
  AL_MUX \picorv32_core/sel15_b12  (
    .i0(\picorv32_core/reg_next_pc [12]),
    .i1(\picorv32_core/n453 [12]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [12]));
  AL_MUX \picorv32_core/sel15_b13  (
    .i0(\picorv32_core/reg_next_pc [13]),
    .i1(\picorv32_core/n453 [13]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [13]));
  AL_MUX \picorv32_core/sel15_b14  (
    .i0(\picorv32_core/reg_next_pc [14]),
    .i1(\picorv32_core/n453 [14]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [14]));
  AL_MUX \picorv32_core/sel15_b15  (
    .i0(\picorv32_core/reg_next_pc [15]),
    .i1(\picorv32_core/n453 [15]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [15]));
  AL_MUX \picorv32_core/sel15_b16  (
    .i0(\picorv32_core/reg_next_pc [16]),
    .i1(\picorv32_core/n453 [16]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [16]));
  AL_MUX \picorv32_core/sel15_b17  (
    .i0(\picorv32_core/reg_next_pc [17]),
    .i1(\picorv32_core/n453 [17]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [17]));
  AL_MUX \picorv32_core/sel15_b18  (
    .i0(\picorv32_core/reg_next_pc [18]),
    .i1(\picorv32_core/n453 [18]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [18]));
  AL_MUX \picorv32_core/sel15_b19  (
    .i0(\picorv32_core/reg_next_pc [19]),
    .i1(\picorv32_core/n453 [19]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [19]));
  AL_MUX \picorv32_core/sel15_b2  (
    .i0(\picorv32_core/reg_next_pc [2]),
    .i1(\picorv32_core/n453 [2]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [2]));
  AL_MUX \picorv32_core/sel15_b20  (
    .i0(\picorv32_core/reg_next_pc [20]),
    .i1(\picorv32_core/n453 [20]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [20]));
  AL_MUX \picorv32_core/sel15_b21  (
    .i0(\picorv32_core/reg_next_pc [21]),
    .i1(\picorv32_core/n453 [21]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [21]));
  AL_MUX \picorv32_core/sel15_b22  (
    .i0(\picorv32_core/reg_next_pc [22]),
    .i1(\picorv32_core/n453 [22]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [22]));
  AL_MUX \picorv32_core/sel15_b23  (
    .i0(\picorv32_core/reg_next_pc [23]),
    .i1(\picorv32_core/n453 [23]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [23]));
  AL_MUX \picorv32_core/sel15_b24  (
    .i0(\picorv32_core/reg_next_pc [24]),
    .i1(\picorv32_core/n453 [24]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [24]));
  AL_MUX \picorv32_core/sel15_b25  (
    .i0(\picorv32_core/reg_next_pc [25]),
    .i1(\picorv32_core/n453 [25]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [25]));
  AL_MUX \picorv32_core/sel15_b26  (
    .i0(\picorv32_core/reg_next_pc [26]),
    .i1(\picorv32_core/n453 [26]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [26]));
  AL_MUX \picorv32_core/sel15_b27  (
    .i0(\picorv32_core/reg_next_pc [27]),
    .i1(\picorv32_core/n453 [27]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [27]));
  AL_MUX \picorv32_core/sel15_b28  (
    .i0(\picorv32_core/reg_next_pc [28]),
    .i1(\picorv32_core/n453 [28]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [28]));
  AL_MUX \picorv32_core/sel15_b29  (
    .i0(\picorv32_core/reg_next_pc [29]),
    .i1(\picorv32_core/n453 [29]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [29]));
  AL_MUX \picorv32_core/sel15_b3  (
    .i0(\picorv32_core/reg_next_pc [3]),
    .i1(\picorv32_core/n453 [3]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [3]));
  AL_MUX \picorv32_core/sel15_b30  (
    .i0(\picorv32_core/reg_next_pc [30]),
    .i1(\picorv32_core/n453 [30]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [30]));
  AL_MUX \picorv32_core/sel15_b31  (
    .i0(\picorv32_core/reg_next_pc [31]),
    .i1(\picorv32_core/n453 [31]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [31]));
  AL_MUX \picorv32_core/sel15_b4  (
    .i0(\picorv32_core/reg_next_pc [4]),
    .i1(\picorv32_core/n453 [4]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [4]));
  AL_MUX \picorv32_core/sel15_b5  (
    .i0(\picorv32_core/reg_next_pc [5]),
    .i1(\picorv32_core/n453 [5]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [5]));
  AL_MUX \picorv32_core/sel15_b6  (
    .i0(\picorv32_core/reg_next_pc [6]),
    .i1(\picorv32_core/n453 [6]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [6]));
  AL_MUX \picorv32_core/sel15_b7  (
    .i0(\picorv32_core/reg_next_pc [7]),
    .i1(\picorv32_core/n453 [7]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [7]));
  AL_MUX \picorv32_core/sel15_b8  (
    .i0(\picorv32_core/reg_next_pc [8]),
    .i1(\picorv32_core/n453 [8]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [8]));
  AL_MUX \picorv32_core/sel15_b9  (
    .i0(\picorv32_core/reg_next_pc [9]),
    .i1(\picorv32_core/n453 [9]),
    .sel(\picorv32_core/sel15_b0_sel_is_3_o ),
    .o(\picorv32_core/n500 [9]));
  and \picorv32_core/sel16_b0/and_b0_0  (\picorv32_core/sel16_b0/B0 , \picorv32_core/count_instr [32], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b0/and_b0_1  (\picorv32_core/sel16_b0/B1 , \picorv32_core/count_instr [0], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b0/and_b0_2  (\picorv32_core/sel16_b0/B2 , \picorv32_core/count_cycle [32], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b0/and_b0_3  (\picorv32_core/sel16_b0/B3 , \picorv32_core/count_cycle [0], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b0/or_B0_B1  (\picorv32_core/sel16_b0/or_B0_B1_o , \picorv32_core/sel16_b0/B0 , \picorv32_core/sel16_b0/B1 );
  or \picorv32_core/sel16_b0/or_B2_B3  (\picorv32_core/sel16_b0/or_B2_B3_o , \picorv32_core/sel16_b0/B2 , \picorv32_core/sel16_b0/B3 );
  or \picorv32_core/sel16_b0/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [0], \picorv32_core/sel16_b0/or_B0_B1_o , \picorv32_core/sel16_b0/or_B2_B3_o );
  and \picorv32_core/sel16_b1/and_b0_0  (\picorv32_core/sel16_b1/B0 , \picorv32_core/count_instr [33], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b1/and_b0_1  (\picorv32_core/sel16_b1/B1 , \picorv32_core/count_instr [1], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b1/and_b0_2  (\picorv32_core/sel16_b1/B2 , \picorv32_core/count_cycle [33], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b1/and_b0_3  (\picorv32_core/sel16_b1/B3 , \picorv32_core/count_cycle [1], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b1/or_B0_B1  (\picorv32_core/sel16_b1/or_B0_B1_o , \picorv32_core/sel16_b1/B0 , \picorv32_core/sel16_b1/B1 );
  or \picorv32_core/sel16_b1/or_B2_B3  (\picorv32_core/sel16_b1/or_B2_B3_o , \picorv32_core/sel16_b1/B2 , \picorv32_core/sel16_b1/B3 );
  or \picorv32_core/sel16_b1/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [1], \picorv32_core/sel16_b1/or_B0_B1_o , \picorv32_core/sel16_b1/or_B2_B3_o );
  and \picorv32_core/sel16_b10/and_b0_0  (\picorv32_core/sel16_b10/B0 , \picorv32_core/count_instr [42], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b10/and_b0_1  (\picorv32_core/sel16_b10/B1 , \picorv32_core/count_instr [10], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b10/and_b0_2  (\picorv32_core/sel16_b10/B2 , \picorv32_core/count_cycle [42], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b10/and_b0_3  (\picorv32_core/sel16_b10/B3 , \picorv32_core/count_cycle [10], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b10/or_B0_B1  (\picorv32_core/sel16_b10/or_B0_B1_o , \picorv32_core/sel16_b10/B0 , \picorv32_core/sel16_b10/B1 );
  or \picorv32_core/sel16_b10/or_B2_B3  (\picorv32_core/sel16_b10/or_B2_B3_o , \picorv32_core/sel16_b10/B2 , \picorv32_core/sel16_b10/B3 );
  or \picorv32_core/sel16_b10/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [10], \picorv32_core/sel16_b10/or_B0_B1_o , \picorv32_core/sel16_b10/or_B2_B3_o );
  and \picorv32_core/sel16_b11/and_b0_0  (\picorv32_core/sel16_b11/B0 , \picorv32_core/count_instr [43], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b11/and_b0_1  (\picorv32_core/sel16_b11/B1 , \picorv32_core/count_instr [11], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b11/and_b0_2  (\picorv32_core/sel16_b11/B2 , \picorv32_core/count_cycle [43], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b11/and_b0_3  (\picorv32_core/sel16_b11/B3 , \picorv32_core/count_cycle [11], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b11/or_B0_B1  (\picorv32_core/sel16_b11/or_B0_B1_o , \picorv32_core/sel16_b11/B0 , \picorv32_core/sel16_b11/B1 );
  or \picorv32_core/sel16_b11/or_B2_B3  (\picorv32_core/sel16_b11/or_B2_B3_o , \picorv32_core/sel16_b11/B2 , \picorv32_core/sel16_b11/B3 );
  or \picorv32_core/sel16_b11/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [11], \picorv32_core/sel16_b11/or_B0_B1_o , \picorv32_core/sel16_b11/or_B2_B3_o );
  and \picorv32_core/sel16_b12/and_b0_0  (\picorv32_core/sel16_b12/B0 , \picorv32_core/count_instr [44], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b12/and_b0_1  (\picorv32_core/sel16_b12/B1 , \picorv32_core/count_instr [12], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b12/and_b0_2  (\picorv32_core/sel16_b12/B2 , \picorv32_core/count_cycle [44], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b12/and_b0_3  (\picorv32_core/sel16_b12/B3 , \picorv32_core/count_cycle [12], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b12/or_B0_B1  (\picorv32_core/sel16_b12/or_B0_B1_o , \picorv32_core/sel16_b12/B0 , \picorv32_core/sel16_b12/B1 );
  or \picorv32_core/sel16_b12/or_B2_B3  (\picorv32_core/sel16_b12/or_B2_B3_o , \picorv32_core/sel16_b12/B2 , \picorv32_core/sel16_b12/B3 );
  or \picorv32_core/sel16_b12/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [12], \picorv32_core/sel16_b12/or_B0_B1_o , \picorv32_core/sel16_b12/or_B2_B3_o );
  and \picorv32_core/sel16_b13/and_b0_0  (\picorv32_core/sel16_b13/B0 , \picorv32_core/count_instr [45], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b13/and_b0_1  (\picorv32_core/sel16_b13/B1 , \picorv32_core/count_instr [13], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b13/and_b0_2  (\picorv32_core/sel16_b13/B2 , \picorv32_core/count_cycle [45], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b13/and_b0_3  (\picorv32_core/sel16_b13/B3 , \picorv32_core/count_cycle [13], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b13/or_B0_B1  (\picorv32_core/sel16_b13/or_B0_B1_o , \picorv32_core/sel16_b13/B0 , \picorv32_core/sel16_b13/B1 );
  or \picorv32_core/sel16_b13/or_B2_B3  (\picorv32_core/sel16_b13/or_B2_B3_o , \picorv32_core/sel16_b13/B2 , \picorv32_core/sel16_b13/B3 );
  or \picorv32_core/sel16_b13/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [13], \picorv32_core/sel16_b13/or_B0_B1_o , \picorv32_core/sel16_b13/or_B2_B3_o );
  and \picorv32_core/sel16_b14/and_b0_0  (\picorv32_core/sel16_b14/B0 , \picorv32_core/count_instr [46], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b14/and_b0_1  (\picorv32_core/sel16_b14/B1 , \picorv32_core/count_instr [14], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b14/and_b0_2  (\picorv32_core/sel16_b14/B2 , \picorv32_core/count_cycle [46], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b14/and_b0_3  (\picorv32_core/sel16_b14/B3 , \picorv32_core/count_cycle [14], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b14/or_B0_B1  (\picorv32_core/sel16_b14/or_B0_B1_o , \picorv32_core/sel16_b14/B0 , \picorv32_core/sel16_b14/B1 );
  or \picorv32_core/sel16_b14/or_B2_B3  (\picorv32_core/sel16_b14/or_B2_B3_o , \picorv32_core/sel16_b14/B2 , \picorv32_core/sel16_b14/B3 );
  or \picorv32_core/sel16_b14/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [14], \picorv32_core/sel16_b14/or_B0_B1_o , \picorv32_core/sel16_b14/or_B2_B3_o );
  and \picorv32_core/sel16_b15/and_b0_0  (\picorv32_core/sel16_b15/B0 , \picorv32_core/count_instr [47], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b15/and_b0_1  (\picorv32_core/sel16_b15/B1 , \picorv32_core/count_instr [15], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b15/and_b0_2  (\picorv32_core/sel16_b15/B2 , \picorv32_core/count_cycle [47], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b15/and_b0_3  (\picorv32_core/sel16_b15/B3 , \picorv32_core/count_cycle [15], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b15/or_B0_B1  (\picorv32_core/sel16_b15/or_B0_B1_o , \picorv32_core/sel16_b15/B0 , \picorv32_core/sel16_b15/B1 );
  or \picorv32_core/sel16_b15/or_B2_B3  (\picorv32_core/sel16_b15/or_B2_B3_o , \picorv32_core/sel16_b15/B2 , \picorv32_core/sel16_b15/B3 );
  or \picorv32_core/sel16_b15/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [15], \picorv32_core/sel16_b15/or_B0_B1_o , \picorv32_core/sel16_b15/or_B2_B3_o );
  and \picorv32_core/sel16_b16/and_b0_0  (\picorv32_core/sel16_b16/B0 , \picorv32_core/count_instr [48], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b16/and_b0_1  (\picorv32_core/sel16_b16/B1 , \picorv32_core/count_instr [16], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b16/and_b0_2  (\picorv32_core/sel16_b16/B2 , \picorv32_core/count_cycle [48], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b16/and_b0_3  (\picorv32_core/sel16_b16/B3 , \picorv32_core/count_cycle [16], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b16/or_B0_B1  (\picorv32_core/sel16_b16/or_B0_B1_o , \picorv32_core/sel16_b16/B0 , \picorv32_core/sel16_b16/B1 );
  or \picorv32_core/sel16_b16/or_B2_B3  (\picorv32_core/sel16_b16/or_B2_B3_o , \picorv32_core/sel16_b16/B2 , \picorv32_core/sel16_b16/B3 );
  or \picorv32_core/sel16_b16/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [16], \picorv32_core/sel16_b16/or_B0_B1_o , \picorv32_core/sel16_b16/or_B2_B3_o );
  and \picorv32_core/sel16_b17/and_b0_0  (\picorv32_core/sel16_b17/B0 , \picorv32_core/count_instr [49], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b17/and_b0_1  (\picorv32_core/sel16_b17/B1 , \picorv32_core/count_instr [17], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b17/and_b0_2  (\picorv32_core/sel16_b17/B2 , \picorv32_core/count_cycle [49], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b17/and_b0_3  (\picorv32_core/sel16_b17/B3 , \picorv32_core/count_cycle [17], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b17/or_B0_B1  (\picorv32_core/sel16_b17/or_B0_B1_o , \picorv32_core/sel16_b17/B0 , \picorv32_core/sel16_b17/B1 );
  or \picorv32_core/sel16_b17/or_B2_B3  (\picorv32_core/sel16_b17/or_B2_B3_o , \picorv32_core/sel16_b17/B2 , \picorv32_core/sel16_b17/B3 );
  or \picorv32_core/sel16_b17/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [17], \picorv32_core/sel16_b17/or_B0_B1_o , \picorv32_core/sel16_b17/or_B2_B3_o );
  and \picorv32_core/sel16_b18/and_b0_0  (\picorv32_core/sel16_b18/B0 , \picorv32_core/count_instr [50], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b18/and_b0_1  (\picorv32_core/sel16_b18/B1 , \picorv32_core/count_instr [18], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b18/and_b0_2  (\picorv32_core/sel16_b18/B2 , \picorv32_core/count_cycle [50], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b18/and_b0_3  (\picorv32_core/sel16_b18/B3 , \picorv32_core/count_cycle [18], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b18/or_B0_B1  (\picorv32_core/sel16_b18/or_B0_B1_o , \picorv32_core/sel16_b18/B0 , \picorv32_core/sel16_b18/B1 );
  or \picorv32_core/sel16_b18/or_B2_B3  (\picorv32_core/sel16_b18/or_B2_B3_o , \picorv32_core/sel16_b18/B2 , \picorv32_core/sel16_b18/B3 );
  or \picorv32_core/sel16_b18/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [18], \picorv32_core/sel16_b18/or_B0_B1_o , \picorv32_core/sel16_b18/or_B2_B3_o );
  and \picorv32_core/sel16_b19/and_b0_0  (\picorv32_core/sel16_b19/B0 , \picorv32_core/count_instr [51], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b19/and_b0_1  (\picorv32_core/sel16_b19/B1 , \picorv32_core/count_instr [19], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b19/and_b0_2  (\picorv32_core/sel16_b19/B2 , \picorv32_core/count_cycle [51], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b19/and_b0_3  (\picorv32_core/sel16_b19/B3 , \picorv32_core/count_cycle [19], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b19/or_B0_B1  (\picorv32_core/sel16_b19/or_B0_B1_o , \picorv32_core/sel16_b19/B0 , \picorv32_core/sel16_b19/B1 );
  or \picorv32_core/sel16_b19/or_B2_B3  (\picorv32_core/sel16_b19/or_B2_B3_o , \picorv32_core/sel16_b19/B2 , \picorv32_core/sel16_b19/B3 );
  or \picorv32_core/sel16_b19/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [19], \picorv32_core/sel16_b19/or_B0_B1_o , \picorv32_core/sel16_b19/or_B2_B3_o );
  and \picorv32_core/sel16_b2/and_b0_0  (\picorv32_core/sel16_b2/B0 , \picorv32_core/count_instr [34], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b2/and_b0_1  (\picorv32_core/sel16_b2/B1 , \picorv32_core/count_instr [2], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b2/and_b0_2  (\picorv32_core/sel16_b2/B2 , \picorv32_core/count_cycle [34], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b2/and_b0_3  (\picorv32_core/sel16_b2/B3 , \picorv32_core/count_cycle [2], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b2/or_B0_B1  (\picorv32_core/sel16_b2/or_B0_B1_o , \picorv32_core/sel16_b2/B0 , \picorv32_core/sel16_b2/B1 );
  or \picorv32_core/sel16_b2/or_B2_B3  (\picorv32_core/sel16_b2/or_B2_B3_o , \picorv32_core/sel16_b2/B2 , \picorv32_core/sel16_b2/B3 );
  or \picorv32_core/sel16_b2/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [2], \picorv32_core/sel16_b2/or_B0_B1_o , \picorv32_core/sel16_b2/or_B2_B3_o );
  and \picorv32_core/sel16_b20/and_b0_0  (\picorv32_core/sel16_b20/B0 , \picorv32_core/count_instr [52], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b20/and_b0_1  (\picorv32_core/sel16_b20/B1 , \picorv32_core/count_instr [20], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b20/and_b0_2  (\picorv32_core/sel16_b20/B2 , \picorv32_core/count_cycle [52], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b20/and_b0_3  (\picorv32_core/sel16_b20/B3 , \picorv32_core/count_cycle [20], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b20/or_B0_B1  (\picorv32_core/sel16_b20/or_B0_B1_o , \picorv32_core/sel16_b20/B0 , \picorv32_core/sel16_b20/B1 );
  or \picorv32_core/sel16_b20/or_B2_B3  (\picorv32_core/sel16_b20/or_B2_B3_o , \picorv32_core/sel16_b20/B2 , \picorv32_core/sel16_b20/B3 );
  or \picorv32_core/sel16_b20/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [20], \picorv32_core/sel16_b20/or_B0_B1_o , \picorv32_core/sel16_b20/or_B2_B3_o );
  and \picorv32_core/sel16_b21/and_b0_0  (\picorv32_core/sel16_b21/B0 , \picorv32_core/count_instr [53], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b21/and_b0_1  (\picorv32_core/sel16_b21/B1 , \picorv32_core/count_instr [21], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b21/and_b0_2  (\picorv32_core/sel16_b21/B2 , \picorv32_core/count_cycle [53], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b21/and_b0_3  (\picorv32_core/sel16_b21/B3 , \picorv32_core/count_cycle [21], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b21/or_B0_B1  (\picorv32_core/sel16_b21/or_B0_B1_o , \picorv32_core/sel16_b21/B0 , \picorv32_core/sel16_b21/B1 );
  or \picorv32_core/sel16_b21/or_B2_B3  (\picorv32_core/sel16_b21/or_B2_B3_o , \picorv32_core/sel16_b21/B2 , \picorv32_core/sel16_b21/B3 );
  or \picorv32_core/sel16_b21/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [21], \picorv32_core/sel16_b21/or_B0_B1_o , \picorv32_core/sel16_b21/or_B2_B3_o );
  and \picorv32_core/sel16_b22/and_b0_0  (\picorv32_core/sel16_b22/B0 , \picorv32_core/count_instr [54], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b22/and_b0_1  (\picorv32_core/sel16_b22/B1 , \picorv32_core/count_instr [22], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b22/and_b0_2  (\picorv32_core/sel16_b22/B2 , \picorv32_core/count_cycle [54], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b22/and_b0_3  (\picorv32_core/sel16_b22/B3 , \picorv32_core/count_cycle [22], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b22/or_B0_B1  (\picorv32_core/sel16_b22/or_B0_B1_o , \picorv32_core/sel16_b22/B0 , \picorv32_core/sel16_b22/B1 );
  or \picorv32_core/sel16_b22/or_B2_B3  (\picorv32_core/sel16_b22/or_B2_B3_o , \picorv32_core/sel16_b22/B2 , \picorv32_core/sel16_b22/B3 );
  or \picorv32_core/sel16_b22/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [22], \picorv32_core/sel16_b22/or_B0_B1_o , \picorv32_core/sel16_b22/or_B2_B3_o );
  and \picorv32_core/sel16_b23/and_b0_0  (\picorv32_core/sel16_b23/B0 , \picorv32_core/count_instr [55], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b23/and_b0_1  (\picorv32_core/sel16_b23/B1 , \picorv32_core/count_instr [23], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b23/and_b0_2  (\picorv32_core/sel16_b23/B2 , \picorv32_core/count_cycle [55], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b23/and_b0_3  (\picorv32_core/sel16_b23/B3 , \picorv32_core/count_cycle [23], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b23/or_B0_B1  (\picorv32_core/sel16_b23/or_B0_B1_o , \picorv32_core/sel16_b23/B0 , \picorv32_core/sel16_b23/B1 );
  or \picorv32_core/sel16_b23/or_B2_B3  (\picorv32_core/sel16_b23/or_B2_B3_o , \picorv32_core/sel16_b23/B2 , \picorv32_core/sel16_b23/B3 );
  or \picorv32_core/sel16_b23/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [23], \picorv32_core/sel16_b23/or_B0_B1_o , \picorv32_core/sel16_b23/or_B2_B3_o );
  and \picorv32_core/sel16_b24/and_b0_0  (\picorv32_core/sel16_b24/B0 , \picorv32_core/count_instr [56], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b24/and_b0_1  (\picorv32_core/sel16_b24/B1 , \picorv32_core/count_instr [24], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b24/and_b0_2  (\picorv32_core/sel16_b24/B2 , \picorv32_core/count_cycle [56], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b24/and_b0_3  (\picorv32_core/sel16_b24/B3 , \picorv32_core/count_cycle [24], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b24/or_B0_B1  (\picorv32_core/sel16_b24/or_B0_B1_o , \picorv32_core/sel16_b24/B0 , \picorv32_core/sel16_b24/B1 );
  or \picorv32_core/sel16_b24/or_B2_B3  (\picorv32_core/sel16_b24/or_B2_B3_o , \picorv32_core/sel16_b24/B2 , \picorv32_core/sel16_b24/B3 );
  or \picorv32_core/sel16_b24/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [24], \picorv32_core/sel16_b24/or_B0_B1_o , \picorv32_core/sel16_b24/or_B2_B3_o );
  and \picorv32_core/sel16_b25/and_b0_0  (\picorv32_core/sel16_b25/B0 , \picorv32_core/count_instr [57], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b25/and_b0_1  (\picorv32_core/sel16_b25/B1 , \picorv32_core/count_instr [25], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b25/and_b0_2  (\picorv32_core/sel16_b25/B2 , \picorv32_core/count_cycle [57], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b25/and_b0_3  (\picorv32_core/sel16_b25/B3 , \picorv32_core/count_cycle [25], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b25/or_B0_B1  (\picorv32_core/sel16_b25/or_B0_B1_o , \picorv32_core/sel16_b25/B0 , \picorv32_core/sel16_b25/B1 );
  or \picorv32_core/sel16_b25/or_B2_B3  (\picorv32_core/sel16_b25/or_B2_B3_o , \picorv32_core/sel16_b25/B2 , \picorv32_core/sel16_b25/B3 );
  or \picorv32_core/sel16_b25/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [25], \picorv32_core/sel16_b25/or_B0_B1_o , \picorv32_core/sel16_b25/or_B2_B3_o );
  and \picorv32_core/sel16_b26/and_b0_0  (\picorv32_core/sel16_b26/B0 , \picorv32_core/count_instr [58], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b26/and_b0_1  (\picorv32_core/sel16_b26/B1 , \picorv32_core/count_instr [26], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b26/and_b0_2  (\picorv32_core/sel16_b26/B2 , \picorv32_core/count_cycle [58], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b26/and_b0_3  (\picorv32_core/sel16_b26/B3 , \picorv32_core/count_cycle [26], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b26/or_B0_B1  (\picorv32_core/sel16_b26/or_B0_B1_o , \picorv32_core/sel16_b26/B0 , \picorv32_core/sel16_b26/B1 );
  or \picorv32_core/sel16_b26/or_B2_B3  (\picorv32_core/sel16_b26/or_B2_B3_o , \picorv32_core/sel16_b26/B2 , \picorv32_core/sel16_b26/B3 );
  or \picorv32_core/sel16_b26/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [26], \picorv32_core/sel16_b26/or_B0_B1_o , \picorv32_core/sel16_b26/or_B2_B3_o );
  and \picorv32_core/sel16_b27/and_b0_0  (\picorv32_core/sel16_b27/B0 , \picorv32_core/count_instr [59], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b27/and_b0_1  (\picorv32_core/sel16_b27/B1 , \picorv32_core/count_instr [27], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b27/and_b0_2  (\picorv32_core/sel16_b27/B2 , \picorv32_core/count_cycle [59], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b27/and_b0_3  (\picorv32_core/sel16_b27/B3 , \picorv32_core/count_cycle [27], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b27/or_B0_B1  (\picorv32_core/sel16_b27/or_B0_B1_o , \picorv32_core/sel16_b27/B0 , \picorv32_core/sel16_b27/B1 );
  or \picorv32_core/sel16_b27/or_B2_B3  (\picorv32_core/sel16_b27/or_B2_B3_o , \picorv32_core/sel16_b27/B2 , \picorv32_core/sel16_b27/B3 );
  or \picorv32_core/sel16_b27/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [27], \picorv32_core/sel16_b27/or_B0_B1_o , \picorv32_core/sel16_b27/or_B2_B3_o );
  and \picorv32_core/sel16_b28/and_b0_0  (\picorv32_core/sel16_b28/B0 , \picorv32_core/count_instr [60], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b28/and_b0_1  (\picorv32_core/sel16_b28/B1 , \picorv32_core/count_instr [28], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b28/and_b0_2  (\picorv32_core/sel16_b28/B2 , \picorv32_core/count_cycle [60], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b28/and_b0_3  (\picorv32_core/sel16_b28/B3 , \picorv32_core/count_cycle [28], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b28/or_B0_B1  (\picorv32_core/sel16_b28/or_B0_B1_o , \picorv32_core/sel16_b28/B0 , \picorv32_core/sel16_b28/B1 );
  or \picorv32_core/sel16_b28/or_B2_B3  (\picorv32_core/sel16_b28/or_B2_B3_o , \picorv32_core/sel16_b28/B2 , \picorv32_core/sel16_b28/B3 );
  or \picorv32_core/sel16_b28/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [28], \picorv32_core/sel16_b28/or_B0_B1_o , \picorv32_core/sel16_b28/or_B2_B3_o );
  and \picorv32_core/sel16_b29/and_b0_0  (\picorv32_core/sel16_b29/B0 , \picorv32_core/count_instr [61], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b29/and_b0_1  (\picorv32_core/sel16_b29/B1 , \picorv32_core/count_instr [29], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b29/and_b0_2  (\picorv32_core/sel16_b29/B2 , \picorv32_core/count_cycle [61], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b29/and_b0_3  (\picorv32_core/sel16_b29/B3 , \picorv32_core/count_cycle [29], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b29/or_B0_B1  (\picorv32_core/sel16_b29/or_B0_B1_o , \picorv32_core/sel16_b29/B0 , \picorv32_core/sel16_b29/B1 );
  or \picorv32_core/sel16_b29/or_B2_B3  (\picorv32_core/sel16_b29/or_B2_B3_o , \picorv32_core/sel16_b29/B2 , \picorv32_core/sel16_b29/B3 );
  or \picorv32_core/sel16_b29/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [29], \picorv32_core/sel16_b29/or_B0_B1_o , \picorv32_core/sel16_b29/or_B2_B3_o );
  and \picorv32_core/sel16_b3/and_b0_0  (\picorv32_core/sel16_b3/B0 , \picorv32_core/count_instr [35], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b3/and_b0_1  (\picorv32_core/sel16_b3/B1 , \picorv32_core/count_instr [3], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b3/and_b0_2  (\picorv32_core/sel16_b3/B2 , \picorv32_core/count_cycle [35], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b3/and_b0_3  (\picorv32_core/sel16_b3/B3 , \picorv32_core/count_cycle [3], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b3/or_B0_B1  (\picorv32_core/sel16_b3/or_B0_B1_o , \picorv32_core/sel16_b3/B0 , \picorv32_core/sel16_b3/B1 );
  or \picorv32_core/sel16_b3/or_B2_B3  (\picorv32_core/sel16_b3/or_B2_B3_o , \picorv32_core/sel16_b3/B2 , \picorv32_core/sel16_b3/B3 );
  or \picorv32_core/sel16_b3/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [3], \picorv32_core/sel16_b3/or_B0_B1_o , \picorv32_core/sel16_b3/or_B2_B3_o );
  and \picorv32_core/sel16_b30/and_b0_0  (\picorv32_core/sel16_b30/B0 , \picorv32_core/count_instr [62], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b30/and_b0_1  (\picorv32_core/sel16_b30/B1 , \picorv32_core/count_instr [30], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b30/and_b0_2  (\picorv32_core/sel16_b30/B2 , \picorv32_core/count_cycle [62], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b30/and_b0_3  (\picorv32_core/sel16_b30/B3 , \picorv32_core/count_cycle [30], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b30/or_B0_B1  (\picorv32_core/sel16_b30/or_B0_B1_o , \picorv32_core/sel16_b30/B0 , \picorv32_core/sel16_b30/B1 );
  or \picorv32_core/sel16_b30/or_B2_B3  (\picorv32_core/sel16_b30/or_B2_B3_o , \picorv32_core/sel16_b30/B2 , \picorv32_core/sel16_b30/B3 );
  or \picorv32_core/sel16_b30/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [30], \picorv32_core/sel16_b30/or_B0_B1_o , \picorv32_core/sel16_b30/or_B2_B3_o );
  and \picorv32_core/sel16_b31/and_b0_0  (\picorv32_core/sel16_b31/B0 , \picorv32_core/count_instr [63], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b31/and_b0_1  (\picorv32_core/sel16_b31/B1 , \picorv32_core/count_instr [31], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b31/and_b0_2  (\picorv32_core/sel16_b31/B2 , \picorv32_core/count_cycle [63], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b31/and_b0_3  (\picorv32_core/sel16_b31/B3 , \picorv32_core/count_cycle [31], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b31/or_B0_B1  (\picorv32_core/sel16_b31/or_B0_B1_o , \picorv32_core/sel16_b31/B0 , \picorv32_core/sel16_b31/B1 );
  or \picorv32_core/sel16_b31/or_B2_B3  (\picorv32_core/sel16_b31/or_B2_B3_o , \picorv32_core/sel16_b31/B2 , \picorv32_core/sel16_b31/B3 );
  or \picorv32_core/sel16_b31/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [31], \picorv32_core/sel16_b31/or_B0_B1_o , \picorv32_core/sel16_b31/or_B2_B3_o );
  and \picorv32_core/sel16_b4/and_b0_0  (\picorv32_core/sel16_b4/B0 , \picorv32_core/count_instr [36], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b4/and_b0_1  (\picorv32_core/sel16_b4/B1 , \picorv32_core/count_instr [4], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b4/and_b0_2  (\picorv32_core/sel16_b4/B2 , \picorv32_core/count_cycle [36], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b4/and_b0_3  (\picorv32_core/sel16_b4/B3 , \picorv32_core/count_cycle [4], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b4/or_B0_B1  (\picorv32_core/sel16_b4/or_B0_B1_o , \picorv32_core/sel16_b4/B0 , \picorv32_core/sel16_b4/B1 );
  or \picorv32_core/sel16_b4/or_B2_B3  (\picorv32_core/sel16_b4/or_B2_B3_o , \picorv32_core/sel16_b4/B2 , \picorv32_core/sel16_b4/B3 );
  or \picorv32_core/sel16_b4/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [4], \picorv32_core/sel16_b4/or_B0_B1_o , \picorv32_core/sel16_b4/or_B2_B3_o );
  and \picorv32_core/sel16_b5/and_b0_0  (\picorv32_core/sel16_b5/B0 , \picorv32_core/count_instr [37], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b5/and_b0_1  (\picorv32_core/sel16_b5/B1 , \picorv32_core/count_instr [5], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b5/and_b0_2  (\picorv32_core/sel16_b5/B2 , \picorv32_core/count_cycle [37], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b5/and_b0_3  (\picorv32_core/sel16_b5/B3 , \picorv32_core/count_cycle [5], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b5/or_B0_B1  (\picorv32_core/sel16_b5/or_B0_B1_o , \picorv32_core/sel16_b5/B0 , \picorv32_core/sel16_b5/B1 );
  or \picorv32_core/sel16_b5/or_B2_B3  (\picorv32_core/sel16_b5/or_B2_B3_o , \picorv32_core/sel16_b5/B2 , \picorv32_core/sel16_b5/B3 );
  or \picorv32_core/sel16_b5/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [5], \picorv32_core/sel16_b5/or_B0_B1_o , \picorv32_core/sel16_b5/or_B2_B3_o );
  and \picorv32_core/sel16_b6/and_b0_0  (\picorv32_core/sel16_b6/B0 , \picorv32_core/count_instr [38], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b6/and_b0_1  (\picorv32_core/sel16_b6/B1 , \picorv32_core/count_instr [6], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b6/and_b0_2  (\picorv32_core/sel16_b6/B2 , \picorv32_core/count_cycle [38], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b6/and_b0_3  (\picorv32_core/sel16_b6/B3 , \picorv32_core/count_cycle [6], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b6/or_B0_B1  (\picorv32_core/sel16_b6/or_B0_B1_o , \picorv32_core/sel16_b6/B0 , \picorv32_core/sel16_b6/B1 );
  or \picorv32_core/sel16_b6/or_B2_B3  (\picorv32_core/sel16_b6/or_B2_B3_o , \picorv32_core/sel16_b6/B2 , \picorv32_core/sel16_b6/B3 );
  or \picorv32_core/sel16_b6/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [6], \picorv32_core/sel16_b6/or_B0_B1_o , \picorv32_core/sel16_b6/or_B2_B3_o );
  and \picorv32_core/sel16_b7/and_b0_0  (\picorv32_core/sel16_b7/B0 , \picorv32_core/count_instr [39], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b7/and_b0_1  (\picorv32_core/sel16_b7/B1 , \picorv32_core/count_instr [7], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b7/and_b0_2  (\picorv32_core/sel16_b7/B2 , \picorv32_core/count_cycle [39], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b7/and_b0_3  (\picorv32_core/sel16_b7/B3 , \picorv32_core/count_cycle [7], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b7/or_B0_B1  (\picorv32_core/sel16_b7/or_B0_B1_o , \picorv32_core/sel16_b7/B0 , \picorv32_core/sel16_b7/B1 );
  or \picorv32_core/sel16_b7/or_B2_B3  (\picorv32_core/sel16_b7/or_B2_B3_o , \picorv32_core/sel16_b7/B2 , \picorv32_core/sel16_b7/B3 );
  or \picorv32_core/sel16_b7/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [7], \picorv32_core/sel16_b7/or_B0_B1_o , \picorv32_core/sel16_b7/or_B2_B3_o );
  and \picorv32_core/sel16_b8/and_b0_0  (\picorv32_core/sel16_b8/B0 , \picorv32_core/count_instr [40], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b8/and_b0_1  (\picorv32_core/sel16_b8/B1 , \picorv32_core/count_instr [8], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b8/and_b0_2  (\picorv32_core/sel16_b8/B2 , \picorv32_core/count_cycle [40], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b8/and_b0_3  (\picorv32_core/sel16_b8/B3 , \picorv32_core/count_cycle [8], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b8/or_B0_B1  (\picorv32_core/sel16_b8/or_B0_B1_o , \picorv32_core/sel16_b8/B0 , \picorv32_core/sel16_b8/B1 );
  or \picorv32_core/sel16_b8/or_B2_B3  (\picorv32_core/sel16_b8/or_B2_B3_o , \picorv32_core/sel16_b8/B2 , \picorv32_core/sel16_b8/B3 );
  or \picorv32_core/sel16_b8/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [8], \picorv32_core/sel16_b8/or_B0_B1_o , \picorv32_core/sel16_b8/or_B2_B3_o );
  and \picorv32_core/sel16_b9/and_b0_0  (\picorv32_core/sel16_b9/B0 , \picorv32_core/count_instr [41], \picorv32_core/instr_rdinstrh );
  and \picorv32_core/sel16_b9/and_b0_1  (\picorv32_core/sel16_b9/B1 , \picorv32_core/count_instr [9], \picorv32_core/instr_rdinstr );
  and \picorv32_core/sel16_b9/and_b0_2  (\picorv32_core/sel16_b9/B2 , \picorv32_core/count_cycle [41], \picorv32_core/instr_rdcycleh );
  and \picorv32_core/sel16_b9/and_b0_3  (\picorv32_core/sel16_b9/B3 , \picorv32_core/count_cycle [9], \picorv32_core/instr_rdcycle );
  or \picorv32_core/sel16_b9/or_B0_B1  (\picorv32_core/sel16_b9/or_B0_B1_o , \picorv32_core/sel16_b9/B0 , \picorv32_core/sel16_b9/B1 );
  or \picorv32_core/sel16_b9/or_B2_B3  (\picorv32_core/sel16_b9/or_B2_B3_o , \picorv32_core/sel16_b9/B2 , \picorv32_core/sel16_b9/B3 );
  or \picorv32_core/sel16_b9/or_or_B0_B1_o_or_B2_  (\picorv32_core/n525 [9], \picorv32_core/sel16_b9/or_B0_B1_o , \picorv32_core/sel16_b9/or_B2_B3_o );
  AL_MUX \picorv32_core/sel17_b1  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\picorv32_core/is_sb_sh_sw ),
    .o(\picorv32_core/n521 [1]));  // ../src/picorv32.v(1690)
  AL_MUX \picorv32_core/sel17_b2  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\picorv32_core/is_sll_srl_sra ),
    .o(\picorv32_core/n521 [2]));  // ../src/picorv32.v(1690)
  AL_MUX \picorv32_core/sel17_b3  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\picorv32_core/n520 ),
    .o(\picorv32_core/n521 [3]));  // ../src/picorv32.v(1690)
  and \picorv32_core/sel18/and_b0_0  (\picorv32_core/sel18/B0 , \picorv32_core/mem_do_prefetch , \picorv32_core/n520 );
  and \picorv32_core/sel18/and_b0_1  (\picorv32_core/sel18/B1 , \picorv32_core/mem_do_rinst , \picorv32_core/is_sll_srl_sra );
  or \picorv32_core/sel18/or_B0_or_B1_B2_o  (\picorv32_core/n522 , \picorv32_core/sel18/B0 , \picorv32_core/sel18/or_B1_B2_o );
  or \picorv32_core/sel18/or_B1_B2  (\picorv32_core/sel18/or_B1_B2_o , \picorv32_core/sel18/B1 , \picorv32_core/is_sb_sh_sw );
  AL_MUX \picorv32_core/sel19_b0  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\picorv32_core/n519 ),
    .o(\picorv32_core/n524 [0]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel19_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/n521 [1]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n524 [1]));  // ../src/picorv32.v(1694)
  and \picorv32_core/sel19_b2/and_b0_0  (\picorv32_core/sel19_b2/B0 , \picorv32_core/n521 [2], \picorv32_core/n523 );
  or \picorv32_core/sel19_b2/or_B0_or_B1_B2_o  (\picorv32_core/sel19_b2/or_B0_or_B1_B2_o_o , \picorv32_core/sel19_b2/B0 , \picorv32_core/is_slli_srli_srai );
  and \picorv32_core/sel19_b3/and_b0_0  (\picorv32_core/sel19_b3/B0 , \picorv32_core/n521 [3], \picorv32_core/n523 );
  or \picorv32_core/sel19_b3/or_B0_or_B1_B2_o  (\picorv32_core/sel19_b3/or_B0_or_B1_B2_o_o , \picorv32_core/sel19_b3/B0 , \picorv32_core/is_jalr_addi_slti_sltiu_xori_ori_andi );
  or \picorv32_core/sel19_b3/or_or_B0_or_B1_B2_o_  (\picorv32_core/n524 [3], \picorv32_core/sel19_b3/or_B0_or_B1_B2_o_o , \picorv32_core/is_lui_auipc_jal );
  AL_MUX \picorv32_core/sel19_b6  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\picorv32_core/is_rdcycle_rdcycleh_rdinstr_rdinstrh ),
    .o(\picorv32_core/n524 [6]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel19_b7  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\picorv32_core/instr_trap ),
    .o(\picorv32_core/n524 [7]));  // ../src/picorv32.v(1694)
  and \picorv32_core/sel1_b0/and_b0_0  (\picorv32_core/sel1_b0/B0 , \picorv32_core/n42 [14], \picorv32_core/n100 );
  and \picorv32_core/sel1_b0/and_b0_1  (\picorv32_core/sel1_b0/B1 , \picorv32_core/n93 [0], \picorv32_core/n98 );
  or \picorv32_core/sel1_b0/or_B0_or_B1_B2_o  (\picorv32_core/n102 [0], \picorv32_core/sel1_b0/B0 , \picorv32_core/sel1_b0/B1 );
  and \picorv32_core/sel1_b1/and_b0_0  (\picorv32_core/sel1_b1/B0 , \picorv32_core/n42 [28], \picorv32_core/n100 );
  and \picorv32_core/sel1_b1/and_b0_1  (\picorv32_core/sel1_b1/B1 , \picorv32_core/n93 [1], \picorv32_core/n98 );
  or \picorv32_core/sel1_b1/or_B0_or_B1_B2_o  (\picorv32_core/n102 [1], \picorv32_core/sel1_b1/B0 , \picorv32_core/sel1_b1/B1 );
  and \picorv32_core/sel1_b2/and_b0_0  (\picorv32_core/sel1_b2/B0 , \picorv32_core/n42 [29], \picorv32_core/n100 );
  and \picorv32_core/sel1_b2/and_b0_1  (\picorv32_core/sel1_b2/B1 , \picorv32_core/n93 [2], \picorv32_core/n98 );
  or \picorv32_core/sel1_b2/or_B0_or_B1_B2_o  (\picorv32_core/n102 [2], \picorv32_core/sel1_b2/B0 , \picorv32_core/sel1_b2/B1 );
  and \picorv32_core/sel1_b3/and_b0_0  (\picorv32_core/sel1_b3/B0 , \picorv32_core/n42 [30], \picorv32_core/n100 );
  and \picorv32_core/sel1_b3/and_b0_1  (\picorv32_core/sel1_b3/B1 , \picorv32_core/n93 [3], \picorv32_core/n98 );
  or \picorv32_core/sel1_b3/or_B0_or_B1_B2_o  (\picorv32_core/n102 [3], \picorv32_core/sel1_b3/B0 , \picorv32_core/sel1_b3/B1 );
  and \picorv32_core/sel1_b4/and_b0_0  (\picorv32_core/sel1_b4/B0 , \picorv32_core/n42 [31], \picorv32_core/n100 );
  and \picorv32_core/sel1_b4/and_b0_1  (\picorv32_core/sel1_b4/B1 , \picorv32_core/n93 [4], \picorv32_core/n98 );
  or \picorv32_core/sel1_b4/or_B0_or_B1_B2_o  (\picorv32_core/n102 [4], \picorv32_core/sel1_b4/B0 , \picorv32_core/sel1_b4/B1 );
  and \picorv32_core/sel2/and_b0_0  (\picorv32_core/sel2/B0 , \picorv32_core/n42 [23], \picorv32_core/n50 );
  and \picorv32_core/sel2/and_b0_1  (\picorv32_core/sel2/B1 , \picorv32_core/mem_rdata_latched [10], \picorv32_core/n97 );
  and \picorv32_core/sel2/and_b0_2  (\picorv32_core/sel2/B2 , \picorv32_core/mem_rdata_latched [5], \picorv32_core/n96 );
  or \picorv32_core/sel2/or_B0_or_B1_B2_o  (\picorv32_core/n51 , \picorv32_core/sel2/B0 , \picorv32_core/sel2/or_B1_B2_o );
  or \picorv32_core/sel2/or_B1_B2  (\picorv32_core/sel2/or_B1_B2_o , \picorv32_core/sel2/B1 , \picorv32_core/sel2/B2 );
  AL_MUX \picorv32_core/sel21_b0  (
    .i0(\picorv32_core/cpuregs_rs1 [0]),
    .i1(\picorv32_core/n518 [0]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [0]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b1  (
    .i0(\picorv32_core/cpuregs_rs1 [1]),
    .i1(\picorv32_core/n518 [1]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [1]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b10  (
    .i0(\picorv32_core/cpuregs_rs1 [10]),
    .i1(\picorv32_core/n518 [10]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [10]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b11  (
    .i0(\picorv32_core/cpuregs_rs1 [11]),
    .i1(\picorv32_core/n518 [11]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [11]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b12  (
    .i0(\picorv32_core/cpuregs_rs1 [12]),
    .i1(\picorv32_core/n518 [12]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [12]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b13  (
    .i0(\picorv32_core/cpuregs_rs1 [13]),
    .i1(\picorv32_core/n518 [13]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [13]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b14  (
    .i0(\picorv32_core/cpuregs_rs1 [14]),
    .i1(\picorv32_core/n518 [14]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [14]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b15  (
    .i0(\picorv32_core/cpuregs_rs1 [15]),
    .i1(\picorv32_core/n518 [15]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [15]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b16  (
    .i0(\picorv32_core/cpuregs_rs1 [16]),
    .i1(\picorv32_core/n518 [16]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [16]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b17  (
    .i0(\picorv32_core/cpuregs_rs1 [17]),
    .i1(\picorv32_core/n518 [17]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [17]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b18  (
    .i0(\picorv32_core/cpuregs_rs1 [18]),
    .i1(\picorv32_core/n518 [18]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [18]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b19  (
    .i0(\picorv32_core/cpuregs_rs1 [19]),
    .i1(\picorv32_core/n518 [19]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [19]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b2  (
    .i0(\picorv32_core/cpuregs_rs1 [2]),
    .i1(\picorv32_core/n518 [2]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [2]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b20  (
    .i0(\picorv32_core/cpuregs_rs1 [20]),
    .i1(\picorv32_core/n518 [20]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [20]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b21  (
    .i0(\picorv32_core/cpuregs_rs1 [21]),
    .i1(\picorv32_core/n518 [21]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [21]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b22  (
    .i0(\picorv32_core/cpuregs_rs1 [22]),
    .i1(\picorv32_core/n518 [22]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [22]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b23  (
    .i0(\picorv32_core/cpuregs_rs1 [23]),
    .i1(\picorv32_core/n518 [23]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [23]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b24  (
    .i0(\picorv32_core/cpuregs_rs1 [24]),
    .i1(\picorv32_core/n518 [24]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [24]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b25  (
    .i0(\picorv32_core/cpuregs_rs1 [25]),
    .i1(\picorv32_core/n518 [25]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [25]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b26  (
    .i0(\picorv32_core/cpuregs_rs1 [26]),
    .i1(\picorv32_core/n518 [26]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [26]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b27  (
    .i0(\picorv32_core/cpuregs_rs1 [27]),
    .i1(\picorv32_core/n518 [27]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [27]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b28  (
    .i0(\picorv32_core/cpuregs_rs1 [28]),
    .i1(\picorv32_core/n518 [28]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [28]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b29  (
    .i0(\picorv32_core/cpuregs_rs1 [29]),
    .i1(\picorv32_core/n518 [29]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [29]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b3  (
    .i0(\picorv32_core/cpuregs_rs1 [3]),
    .i1(\picorv32_core/n518 [3]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [3]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b30  (
    .i0(\picorv32_core/cpuregs_rs1 [30]),
    .i1(\picorv32_core/n518 [30]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [30]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b31  (
    .i0(\picorv32_core/cpuregs_rs1 [31]),
    .i1(\picorv32_core/n518 [31]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [31]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b4  (
    .i0(\picorv32_core/cpuregs_rs1 [4]),
    .i1(\picorv32_core/n518 [4]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [4]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b5  (
    .i0(\picorv32_core/cpuregs_rs1 [5]),
    .i1(\picorv32_core/n518 [5]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [5]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b6  (
    .i0(\picorv32_core/cpuregs_rs1 [6]),
    .i1(\picorv32_core/n518 [6]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [6]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b7  (
    .i0(\picorv32_core/cpuregs_rs1 [7]),
    .i1(\picorv32_core/n518 [7]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [7]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b8  (
    .i0(\picorv32_core/cpuregs_rs1 [8]),
    .i1(\picorv32_core/n518 [8]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [8]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel21_b9  (
    .i0(\picorv32_core/cpuregs_rs1 [9]),
    .i1(\picorv32_core/n518 [9]),
    .sel(\picorv32_core/is_lui_auipc_jal ),
    .o(\picorv32_core/n527 [9]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b0  (
    .i0(\picorv32_core/decoded_imm [0]),
    .i1(\picorv32_core/cpuregs_rs2 [0]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [0]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b1  (
    .i0(\picorv32_core/decoded_imm [1]),
    .i1(\picorv32_core/cpuregs_rs2 [1]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [1]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b10  (
    .i0(\picorv32_core/decoded_imm [10]),
    .i1(\picorv32_core/cpuregs_rs2 [10]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [10]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b11  (
    .i0(\picorv32_core/decoded_imm [11]),
    .i1(\picorv32_core/cpuregs_rs2 [11]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [11]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b12  (
    .i0(\picorv32_core/decoded_imm [12]),
    .i1(\picorv32_core/cpuregs_rs2 [12]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [12]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b13  (
    .i0(\picorv32_core/decoded_imm [13]),
    .i1(\picorv32_core/cpuregs_rs2 [13]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [13]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b14  (
    .i0(\picorv32_core/decoded_imm [14]),
    .i1(\picorv32_core/cpuregs_rs2 [14]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [14]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b15  (
    .i0(\picorv32_core/decoded_imm [15]),
    .i1(\picorv32_core/cpuregs_rs2 [15]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [15]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b16  (
    .i0(\picorv32_core/decoded_imm [16]),
    .i1(\picorv32_core/cpuregs_rs2 [16]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [16]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b17  (
    .i0(\picorv32_core/decoded_imm [17]),
    .i1(\picorv32_core/cpuregs_rs2 [17]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [17]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b18  (
    .i0(\picorv32_core/decoded_imm [18]),
    .i1(\picorv32_core/cpuregs_rs2 [18]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [18]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b19  (
    .i0(\picorv32_core/decoded_imm [19]),
    .i1(\picorv32_core/cpuregs_rs2 [19]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [19]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b2  (
    .i0(\picorv32_core/decoded_imm [2]),
    .i1(\picorv32_core/cpuregs_rs2 [2]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [2]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b20  (
    .i0(\picorv32_core/decoded_imm [20]),
    .i1(\picorv32_core/cpuregs_rs2 [20]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [20]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b21  (
    .i0(\picorv32_core/decoded_imm [21]),
    .i1(\picorv32_core/cpuregs_rs2 [21]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [21]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b22  (
    .i0(\picorv32_core/decoded_imm [22]),
    .i1(\picorv32_core/cpuregs_rs2 [22]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [22]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b23  (
    .i0(\picorv32_core/decoded_imm [23]),
    .i1(\picorv32_core/cpuregs_rs2 [23]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [23]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b24  (
    .i0(\picorv32_core/decoded_imm [24]),
    .i1(\picorv32_core/cpuregs_rs2 [24]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [24]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b25  (
    .i0(\picorv32_core/decoded_imm [25]),
    .i1(\picorv32_core/cpuregs_rs2 [25]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [25]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b26  (
    .i0(\picorv32_core/decoded_imm [26]),
    .i1(\picorv32_core/cpuregs_rs2 [26]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [26]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b27  (
    .i0(\picorv32_core/decoded_imm [27]),
    .i1(\picorv32_core/cpuregs_rs2 [27]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [27]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b28  (
    .i0(\picorv32_core/decoded_imm [28]),
    .i1(\picorv32_core/cpuregs_rs2 [28]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [28]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b29  (
    .i0(\picorv32_core/decoded_imm [29]),
    .i1(\picorv32_core/cpuregs_rs2 [29]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [29]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b3  (
    .i0(\picorv32_core/decoded_imm [3]),
    .i1(\picorv32_core/cpuregs_rs2 [3]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [3]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b30  (
    .i0(\picorv32_core/decoded_imm [30]),
    .i1(\picorv32_core/cpuregs_rs2 [30]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [30]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b31  (
    .i0(\picorv32_core/decoded_imm [31]),
    .i1(\picorv32_core/cpuregs_rs2 [31]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [31]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b4  (
    .i0(\picorv32_core/decoded_imm [4]),
    .i1(\picorv32_core/cpuregs_rs2 [4]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [4]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b5  (
    .i0(\picorv32_core/decoded_imm [5]),
    .i1(\picorv32_core/cpuregs_rs2 [5]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [5]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b6  (
    .i0(\picorv32_core/decoded_imm [6]),
    .i1(\picorv32_core/cpuregs_rs2 [6]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [6]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b7  (
    .i0(\picorv32_core/decoded_imm [7]),
    .i1(\picorv32_core/cpuregs_rs2 [7]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [7]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b8  (
    .i0(\picorv32_core/decoded_imm [8]),
    .i1(\picorv32_core/cpuregs_rs2 [8]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [8]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel22_b9  (
    .i0(\picorv32_core/decoded_imm [9]),
    .i1(\picorv32_core/cpuregs_rs2 [9]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n528 [9]));  // ../src/picorv32.v(1694)
  and \picorv32_core/sel23/and_b0_0  (\picorv32_core/sel23/B0 , \picorv32_core/n522 , \picorv32_core/n523 );
  and \picorv32_core/sel23/and_b0_2  (\picorv32_core/sel23/B2 , \picorv32_core/mem_do_prefetch , \picorv32_core/n530 );
  and \picorv32_core/sel23/and_b0_3  (\picorv32_core/sel23/B3 , \picorv32_core/mem_do_rinst , \picorv32_core/n529 );
  or \picorv32_core/sel23/or_B0_B1  (\picorv32_core/sel23/or_B0_B1_o , \picorv32_core/sel23/B0 , \picorv32_core/n519 );
  or \picorv32_core/sel23/or_B2_B3  (\picorv32_core/sel23/or_B2_B3_o , \picorv32_core/sel23/B2 , \picorv32_core/sel23/B3 );
  or \picorv32_core/sel23/or_or_B0_B1_o_or_B2_  (\picorv32_core/n531 , \picorv32_core/sel23/or_B0_B1_o , \picorv32_core/sel23/or_B2_B3_o );
  AL_MUX \picorv32_core/sel24_b0  (
    .i0(\picorv32_core/decoded_rs2 [0]),
    .i1(\picorv32_core/cpuregs_rs2 [0]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n532 [0]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel24_b1  (
    .i0(\picorv32_core/decoded_rs2 [1]),
    .i1(\picorv32_core/cpuregs_rs2 [1]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n532 [1]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel24_b2  (
    .i0(\picorv32_core/decoded_rs2 [2]),
    .i1(\picorv32_core/cpuregs_rs2 [2]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n532 [2]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel24_b3  (
    .i0(\picorv32_core/decoded_rs2 [3]),
    .i1(\picorv32_core/cpuregs_rs2 [3]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n532 [3]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel24_b4  (
    .i0(\picorv32_core/decoded_rs2 [4]),
    .i1(\picorv32_core/cpuregs_rs2 [4]),
    .sel(\picorv32_core/n523 ),
    .o(\picorv32_core/n532 [4]));  // ../src/picorv32.v(1694)
  AL_MUX \picorv32_core/sel25_b0  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\picorv32_core/instr_sh ),
    .o(\picorv32_core/n575 [0]));  // ../src/picorv32.v(1802)
  AL_MUX \picorv32_core/sel25_b1  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\picorv32_core/instr_sb ),
    .o(\picorv32_core/n575 [1]));  // ../src/picorv32.v(1802)
  AL_MUX \picorv32_core/sel26_b0  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\picorv32_core/n600 ),
    .o(\picorv32_core/n601 [0]));  // ../src/picorv32.v(1827)
  AL_MUX \picorv32_core/sel26_b1  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\picorv32_core/n599 ),
    .o(\picorv32_core/n601 [1]));  // ../src/picorv32.v(1827)
  AL_MUX \picorv32_core/sel27_b10  (
    .i0(\picorv32_core/mem_rdata_word [10]),
    .i1(\picorv32_core/n641 [7]),
    .sel(\picorv32_core/latched_is_lb ),
    .o(\picorv32_core/n641 [10]));  // ../src/picorv32.v(1844)
  AL_MUX \picorv32_core/sel27_b11  (
    .i0(\picorv32_core/mem_rdata_word [11]),
    .i1(\picorv32_core/n641 [7]),
    .sel(\picorv32_core/latched_is_lb ),
    .o(\picorv32_core/n641 [11]));  // ../src/picorv32.v(1844)
  AL_MUX \picorv32_core/sel27_b12  (
    .i0(\picorv32_core/mem_rdata_word [12]),
    .i1(\picorv32_core/n641 [7]),
    .sel(\picorv32_core/latched_is_lb ),
    .o(\picorv32_core/n641 [12]));  // ../src/picorv32.v(1844)
  AL_MUX \picorv32_core/sel27_b13  (
    .i0(\picorv32_core/mem_rdata_word [13]),
    .i1(\picorv32_core/n641 [7]),
    .sel(\picorv32_core/latched_is_lb ),
    .o(\picorv32_core/n641 [13]));  // ../src/picorv32.v(1844)
  AL_MUX \picorv32_core/sel27_b14  (
    .i0(\picorv32_core/mem_rdata_word [14]),
    .i1(\picorv32_core/n641 [7]),
    .sel(\picorv32_core/latched_is_lb ),
    .o(\picorv32_core/n641 [14]));  // ../src/picorv32.v(1844)
  AL_MUX \picorv32_core/sel27_b15  (
    .i0(\picorv32_core/mem_rdata_word [15]),
    .i1(\picorv32_core/n641 [7]),
    .sel(\picorv32_core/latched_is_lb ),
    .o(\picorv32_core/n641 [15]));  // ../src/picorv32.v(1844)
  and \picorv32_core/sel27_b16/and_b0_0  (\picorv32_core/sel27_b16/B0 , \picorv32_core/n641 [7], \picorv32_core/latched_is_lb );
  and \picorv32_core/sel27_b16/and_b0_1  (\picorv32_core/sel27_b16/B1 , \picorv32_core/mem_rdata_word [15], \picorv32_core/latched_is_lh );
  and \picorv32_core/sel27_b16/and_b0_2  (\picorv32_core/sel27_b16/B2 , \picorv32_core/mem_rdata_word [16], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b16/or_B0_or_B1_B2_o  (\picorv32_core/n641 [16], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b16/or_B1_B2_o );
  or \picorv32_core/sel27_b16/or_B1_B2  (\picorv32_core/sel27_b16/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b16/B2 );
  and \picorv32_core/sel27_b17/and_b0_2  (\picorv32_core/sel27_b17/B2 , \picorv32_core/mem_rdata_word [17], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b17/or_B0_or_B1_B2_o  (\picorv32_core/n641 [17], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b17/or_B1_B2_o );
  or \picorv32_core/sel27_b17/or_B1_B2  (\picorv32_core/sel27_b17/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b17/B2 );
  and \picorv32_core/sel27_b18/and_b0_2  (\picorv32_core/sel27_b18/B2 , \picorv32_core/mem_rdata_word [18], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b18/or_B0_or_B1_B2_o  (\picorv32_core/n641 [18], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b18/or_B1_B2_o );
  or \picorv32_core/sel27_b18/or_B1_B2  (\picorv32_core/sel27_b18/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b18/B2 );
  and \picorv32_core/sel27_b19/and_b0_2  (\picorv32_core/sel27_b19/B2 , \picorv32_core/mem_rdata_word [19], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b19/or_B0_or_B1_B2_o  (\picorv32_core/n641 [19], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b19/or_B1_B2_o );
  or \picorv32_core/sel27_b19/or_B1_B2  (\picorv32_core/sel27_b19/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b19/B2 );
  and \picorv32_core/sel27_b20/and_b0_2  (\picorv32_core/sel27_b20/B2 , \picorv32_core/mem_rdata_word [20], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b20/or_B0_or_B1_B2_o  (\picorv32_core/n641 [20], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b20/or_B1_B2_o );
  or \picorv32_core/sel27_b20/or_B1_B2  (\picorv32_core/sel27_b20/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b20/B2 );
  and \picorv32_core/sel27_b21/and_b0_2  (\picorv32_core/sel27_b21/B2 , \picorv32_core/mem_rdata_word [21], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b21/or_B0_or_B1_B2_o  (\picorv32_core/n641 [21], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b21/or_B1_B2_o );
  or \picorv32_core/sel27_b21/or_B1_B2  (\picorv32_core/sel27_b21/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b21/B2 );
  and \picorv32_core/sel27_b22/and_b0_2  (\picorv32_core/sel27_b22/B2 , \picorv32_core/mem_rdata_word [22], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b22/or_B0_or_B1_B2_o  (\picorv32_core/n641 [22], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b22/or_B1_B2_o );
  or \picorv32_core/sel27_b22/or_B1_B2  (\picorv32_core/sel27_b22/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b22/B2 );
  and \picorv32_core/sel27_b23/and_b0_2  (\picorv32_core/sel27_b23/B2 , \picorv32_core/mem_rdata_word [23], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b23/or_B0_or_B1_B2_o  (\picorv32_core/n641 [23], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b23/or_B1_B2_o );
  or \picorv32_core/sel27_b23/or_B1_B2  (\picorv32_core/sel27_b23/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b23/B2 );
  and \picorv32_core/sel27_b24/and_b0_2  (\picorv32_core/sel27_b24/B2 , \picorv32_core/mem_rdata_word [24], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b24/or_B0_or_B1_B2_o  (\picorv32_core/n641 [24], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b24/or_B1_B2_o );
  or \picorv32_core/sel27_b24/or_B1_B2  (\picorv32_core/sel27_b24/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b24/B2 );
  and \picorv32_core/sel27_b25/and_b0_2  (\picorv32_core/sel27_b25/B2 , \picorv32_core/mem_rdata_word [25], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b25/or_B0_or_B1_B2_o  (\picorv32_core/n641 [25], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b25/or_B1_B2_o );
  or \picorv32_core/sel27_b25/or_B1_B2  (\picorv32_core/sel27_b25/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b25/B2 );
  and \picorv32_core/sel27_b26/and_b0_2  (\picorv32_core/sel27_b26/B2 , \picorv32_core/mem_rdata_word [26], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b26/or_B0_or_B1_B2_o  (\picorv32_core/n641 [26], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b26/or_B1_B2_o );
  or \picorv32_core/sel27_b26/or_B1_B2  (\picorv32_core/sel27_b26/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b26/B2 );
  and \picorv32_core/sel27_b27/and_b0_2  (\picorv32_core/sel27_b27/B2 , \picorv32_core/mem_rdata_word [27], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b27/or_B0_or_B1_B2_o  (\picorv32_core/n641 [27], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b27/or_B1_B2_o );
  or \picorv32_core/sel27_b27/or_B1_B2  (\picorv32_core/sel27_b27/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b27/B2 );
  and \picorv32_core/sel27_b28/and_b0_2  (\picorv32_core/sel27_b28/B2 , \picorv32_core/mem_rdata_word [28], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b28/or_B0_or_B1_B2_o  (\picorv32_core/n641 [28], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b28/or_B1_B2_o );
  or \picorv32_core/sel27_b28/or_B1_B2  (\picorv32_core/sel27_b28/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b28/B2 );
  and \picorv32_core/sel27_b29/and_b0_2  (\picorv32_core/sel27_b29/B2 , \picorv32_core/mem_rdata_word [29], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b29/or_B0_or_B1_B2_o  (\picorv32_core/n641 [29], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b29/or_B1_B2_o );
  or \picorv32_core/sel27_b29/or_B1_B2  (\picorv32_core/sel27_b29/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b29/B2 );
  and \picorv32_core/sel27_b30/and_b0_2  (\picorv32_core/sel27_b30/B2 , \picorv32_core/mem_rdata_word [30], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b30/or_B0_or_B1_B2_o  (\picorv32_core/n641 [30], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b30/or_B1_B2_o );
  or \picorv32_core/sel27_b30/or_B1_B2  (\picorv32_core/sel27_b30/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b30/B2 );
  and \picorv32_core/sel27_b31/and_b0_2  (\picorv32_core/sel27_b31/B2 , \picorv32_core/mem_rdata_word [31], \picorv32_core/latched_is_lu );
  or \picorv32_core/sel27_b31/or_B0_or_B1_B2_o  (\picorv32_core/n641 [31], \picorv32_core/sel27_b16/B0 , \picorv32_core/sel27_b31/or_B1_B2_o );
  or \picorv32_core/sel27_b31/or_B1_B2  (\picorv32_core/sel27_b31/or_B1_B2_o , \picorv32_core/sel27_b16/B1 , \picorv32_core/sel27_b31/B2 );
  AL_MUX \picorv32_core/sel27_b8  (
    .i0(\picorv32_core/mem_rdata_word [8]),
    .i1(\picorv32_core/n641 [7]),
    .sel(\picorv32_core/latched_is_lb ),
    .o(\picorv32_core/n641 [8]));  // ../src/picorv32.v(1844)
  AL_MUX \picorv32_core/sel27_b9  (
    .i0(\picorv32_core/mem_rdata_word [9]),
    .i1(\picorv32_core/n641 [7]),
    .sel(\picorv32_core/latched_is_lb ),
    .o(\picorv32_core/n641 [9]));  // ../src/picorv32.v(1844)
  and \picorv32_core/sel28/and_b0_0  (\picorv32_core/sel28/B0 , \picorv32_core/n568 , \picorv32_core/n667 );
  and \picorv32_core/sel28/and_b0_1  (\picorv32_core/sel28/B1 , \picorv32_core/n522 , \picorv32_core/n665 );
  and \picorv32_core/sel28/and_b0_2  (\picorv32_core/sel28/B2 , \picorv32_core/n531 , \picorv32_core/n664 );
  and \picorv32_core/sel28/and_b0_3  (\picorv32_core/sel28/B3 , \picorv32_core/n513 , \picorv32_core/n663 );
  and \picorv32_core/sel28/and_b0_4  (\picorv32_core/sel28/B4 , \picorv32_core/mem_do_rinst , \picorv32_core/n670 );
  or \picorv32_core/sel28/or_B0_B1  (\picorv32_core/sel28/or_B0_B1_o , \picorv32_core/sel28/B0 , \picorv32_core/sel28/B1 );
  or \picorv32_core/sel28/or_B2_or_B3_B4_o  (\picorv32_core/sel28/or_B2_or_B3_B4_o_o , \picorv32_core/sel28/B2 , \picorv32_core/sel28/or_B3_B4_o );
  or \picorv32_core/sel28/or_B3_B4  (\picorv32_core/sel28/or_B3_B4_o , \picorv32_core/sel28/B3 , \picorv32_core/sel28/B4 );
  or \picorv32_core/sel28/or_or_B0_B1_o_or_B2_  (\picorv32_core/n671 , \picorv32_core/sel28/or_B0_B1_o , \picorv32_core/sel28/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel29_b0/and_b0_0  (\picorv32_core/sel29_b0/B0 , \picorv32_core/n652 [0], \picorv32_core/n669 );
  and \picorv32_core/sel29_b0/and_b0_1  (\picorv32_core/sel29_b0/B1 , \picorv32_core/n583 [0], \picorv32_core/n668 );
  and \picorv32_core/sel29_b0/and_b0_2  (\picorv32_core/sel29_b0/B2 , \picorv32_core/mem_wordsize [0], \picorv32_core/n667 );
  and \picorv32_core/sel29_b0/and_b0_3  (\picorv32_core/sel29_b0/B3 , \picorv32_core/mem_wordsize [0], \picorv32_core/n666 );
  and \picorv32_core/sel29_b0/and_b0_4  (\picorv32_core/sel29_b0/B4 , \picorv32_core/mem_wordsize [0], \picorv32_core/n665 );
  and \picorv32_core/sel29_b0/and_b0_5  (\picorv32_core/sel29_b0/B5 , \picorv32_core/mem_wordsize [0], \picorv32_core/n664 );
  and \picorv32_core/sel29_b0/and_b0_7  (\picorv32_core/sel29_b0/B7 , \picorv32_core/mem_wordsize [0], \picorv32_core/n662 );
  or \picorv32_core/sel29_b0/or_B0_B1  (\picorv32_core/sel29_b0/or_B0_B1_o , \picorv32_core/sel29_b0/B0 , \picorv32_core/sel29_b0/B1 );
  or \picorv32_core/sel29_b0/or_B2_B3  (\picorv32_core/sel29_b0/or_B2_B3_o , \picorv32_core/sel29_b0/B2 , \picorv32_core/sel29_b0/B3 );
  or \picorv32_core/sel29_b0/or_B4_B5  (\picorv32_core/sel29_b0/or_B4_B5_o , \picorv32_core/sel29_b0/B4 , \picorv32_core/sel29_b0/B5 );
  or \picorv32_core/sel29_b0/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel29_b0/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel29_b0/or_B0_B1_o , \picorv32_core/sel29_b0/or_B2_B3_o );
  or \picorv32_core/sel29_b0/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel29_b0/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel29_b0/or_B4_B5_o , \picorv32_core/sel29_b0/B7 );
  or \picorv32_core/sel29_b0/or_or_or_B0_B1_o_or_  (\picorv32_core/n672 [0], \picorv32_core/sel29_b0/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel29_b0/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel29_b1/and_b0_0  (\picorv32_core/sel29_b1/B0 , \picorv32_core/n652 [1], \picorv32_core/n669 );
  and \picorv32_core/sel29_b1/and_b0_1  (\picorv32_core/sel29_b1/B1 , \picorv32_core/n583 [1], \picorv32_core/n668 );
  and \picorv32_core/sel29_b1/and_b0_2  (\picorv32_core/sel29_b1/B2 , \picorv32_core/mem_wordsize [1], \picorv32_core/n667 );
  and \picorv32_core/sel29_b1/and_b0_3  (\picorv32_core/sel29_b1/B3 , \picorv32_core/mem_wordsize [1], \picorv32_core/n666 );
  and \picorv32_core/sel29_b1/and_b0_4  (\picorv32_core/sel29_b1/B4 , \picorv32_core/mem_wordsize [1], \picorv32_core/n665 );
  and \picorv32_core/sel29_b1/and_b0_5  (\picorv32_core/sel29_b1/B5 , \picorv32_core/mem_wordsize [1], \picorv32_core/n664 );
  and \picorv32_core/sel29_b1/and_b0_7  (\picorv32_core/sel29_b1/B7 , \picorv32_core/mem_wordsize [1], \picorv32_core/n662 );
  or \picorv32_core/sel29_b1/or_B0_B1  (\picorv32_core/sel29_b1/or_B0_B1_o , \picorv32_core/sel29_b1/B0 , \picorv32_core/sel29_b1/B1 );
  or \picorv32_core/sel29_b1/or_B2_B3  (\picorv32_core/sel29_b1/or_B2_B3_o , \picorv32_core/sel29_b1/B2 , \picorv32_core/sel29_b1/B3 );
  or \picorv32_core/sel29_b1/or_B4_B5  (\picorv32_core/sel29_b1/or_B4_B5_o , \picorv32_core/sel29_b1/B4 , \picorv32_core/sel29_b1/B5 );
  or \picorv32_core/sel29_b1/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel29_b1/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel29_b1/or_B0_B1_o , \picorv32_core/sel29_b1/or_B2_B3_o );
  or \picorv32_core/sel29_b1/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel29_b1/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel29_b1/or_B4_B5_o , \picorv32_core/sel29_b1/B7 );
  or \picorv32_core/sel29_b1/or_or_or_B0_B1_o_or_  (\picorv32_core/n672 [1], \picorv32_core/sel29_b1/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel29_b1/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel32/and_b0_1  (\picorv32_core/sel32/B1 , \picorv32_core/n547 , \picorv32_core/n666 );
  and \picorv32_core/sel32/and_b0_2  (\picorv32_core/sel32/B2 , \picorv32_core/n526 , \picorv32_core/n664 );
  and \picorv32_core/sel32/and_b0_4  (\picorv32_core/sel32/B4 , \picorv32_core/latched_store , \picorv32_core/n675 );
  or \picorv32_core/sel32/or_B0_B1  (\picorv32_core/sel32/or_B0_B1_o , \picorv32_core/n676 , \picorv32_core/sel32/B1 );
  or \picorv32_core/sel32/or_B2_or_B3_B4_o  (\picorv32_core/sel32/or_B2_or_B3_B4_o_o , \picorv32_core/sel32/B2 , \picorv32_core/sel32/B4 );
  or \picorv32_core/sel32/or_or_B0_B1_o_or_B2_  (\picorv32_core/n677 , \picorv32_core/sel32/or_B0_B1_o , \picorv32_core/sel32/or_B2_or_B3_B4_o_o );
  and \picorv32_core/sel33/and_b0_0  (\picorv32_core/sel33/B0 , \picorv32_core/n552 , \picorv32_core/n666 );
  and \picorv32_core/sel33/and_b0_2  (\picorv32_core/sel33/B2 , \picorv32_core/latched_stalu , \picorv32_core/n678 );
  or \picorv32_core/sel33/or_B0_or_B1_B2_o  (\picorv32_core/n679 , \picorv32_core/sel33/B0 , \picorv32_core/sel33/B2 );
  and \picorv32_core/sel34/and_b0_0  (\picorv32_core/sel34/B0 , \picorv32_core/n548 , \picorv32_core/n666 );
  and \picorv32_core/sel34/and_b0_1  (\picorv32_core/sel34/B1 , \picorv32_core/n514 , \picorv32_core/n663 );
  and \picorv32_core/sel34/and_b0_2  (\picorv32_core/sel34/B2 , \picorv32_core/latched_branch , \picorv32_core/n678 );
  or \picorv32_core/sel34/or_B0_or_B1_B2_o  (\picorv32_core/n681 , \picorv32_core/sel34/B0 , \picorv32_core/sel34/or_B1_B2_o );
  or \picorv32_core/sel34/or_B1_B2  (\picorv32_core/sel34/or_B1_B2_o , \picorv32_core/sel34/B1 , \picorv32_core/sel34/B2 );
  and \picorv32_core/sel35/and_b0_0  (\picorv32_core/sel35/B0 , \picorv32_core/n653 , \picorv32_core/n669 );
  and \picorv32_core/sel35/and_b0_2  (\picorv32_core/sel35/B2 , \picorv32_core/latched_is_lu , \picorv32_core/n682 );
  or \picorv32_core/sel35/or_B0_or_B1_B2_o  (\picorv32_core/n683 , \picorv32_core/sel35/B0 , \picorv32_core/sel35/B2 );
  and \picorv32_core/sel36/and_b0_0  (\picorv32_core/sel36/B0 , \picorv32_core/n654 , \picorv32_core/n669 );
  and \picorv32_core/sel36/and_b0_2  (\picorv32_core/sel36/B2 , \picorv32_core/latched_is_lh , \picorv32_core/n682 );
  or \picorv32_core/sel36/or_B0_or_B1_B2_o  (\picorv32_core/n685 , \picorv32_core/sel36/B0 , \picorv32_core/sel36/B2 );
  and \picorv32_core/sel37/and_b0_0  (\picorv32_core/sel37/B0 , \picorv32_core/n655 , \picorv32_core/n669 );
  and \picorv32_core/sel37/and_b0_2  (\picorv32_core/sel37/B2 , \picorv32_core/latched_is_lb , \picorv32_core/n682 );
  or \picorv32_core/sel37/or_B0_or_B1_B2_o  (\picorv32_core/n687 , \picorv32_core/sel37/B0 , \picorv32_core/sel37/B2 );
  and \picorv32_core/sel38_b0/and_b0_0  (\picorv32_core/sel38_b0/B0 , \picorv32_core/latched_rd [0], \picorv32_core/n669 );
  and \picorv32_core/sel38_b0/and_b0_1  (\picorv32_core/sel38_b0/B1 , \picorv32_core/latched_rd [0], \picorv32_core/n668 );
  and \picorv32_core/sel38_b0/and_b0_2  (\picorv32_core/sel38_b0/B2 , \picorv32_core/latched_rd [0], \picorv32_core/n667 );
  and \picorv32_core/sel38_b0/and_b0_3  (\picorv32_core/sel38_b0/B3 , \picorv32_core/n546 [0], \picorv32_core/n666 );
  and \picorv32_core/sel38_b0/and_b0_4  (\picorv32_core/sel38_b0/B4 , \picorv32_core/latched_rd [0], \picorv32_core/n665 );
  and \picorv32_core/sel38_b0/and_b0_5  (\picorv32_core/sel38_b0/B5 , \picorv32_core/latched_rd [0], \picorv32_core/n664 );
  and \picorv32_core/sel38_b0/and_b0_6  (\picorv32_core/sel38_b0/B6 , \picorv32_core/decoded_rd [0], \picorv32_core/n663 );
  and \picorv32_core/sel38_b0/and_b0_7  (\picorv32_core/sel38_b0/B7 , \picorv32_core/latched_rd [0], \picorv32_core/n662 );
  or \picorv32_core/sel38_b0/or_B0_B1  (\picorv32_core/sel38_b0/or_B0_B1_o , \picorv32_core/sel38_b0/B0 , \picorv32_core/sel38_b0/B1 );
  or \picorv32_core/sel38_b0/or_B2_B3  (\picorv32_core/sel38_b0/or_B2_B3_o , \picorv32_core/sel38_b0/B2 , \picorv32_core/sel38_b0/B3 );
  or \picorv32_core/sel38_b0/or_B4_B5  (\picorv32_core/sel38_b0/or_B4_B5_o , \picorv32_core/sel38_b0/B4 , \picorv32_core/sel38_b0/B5 );
  or \picorv32_core/sel38_b0/or_B6_B7  (\picorv32_core/sel38_b0/or_B6_B7_o , \picorv32_core/sel38_b0/B6 , \picorv32_core/sel38_b0/B7 );
  or \picorv32_core/sel38_b0/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel38_b0/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel38_b0/or_B0_B1_o , \picorv32_core/sel38_b0/or_B2_B3_o );
  or \picorv32_core/sel38_b0/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel38_b0/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel38_b0/or_B4_B5_o , \picorv32_core/sel38_b0/or_B6_B7_o );
  or \picorv32_core/sel38_b0/or_or_or_B0_B1_o_or_  (\picorv32_core/n688 [0], \picorv32_core/sel38_b0/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel38_b0/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel38_b1/and_b0_0  (\picorv32_core/sel38_b1/B0 , \picorv32_core/latched_rd [1], \picorv32_core/n669 );
  and \picorv32_core/sel38_b1/and_b0_1  (\picorv32_core/sel38_b1/B1 , \picorv32_core/latched_rd [1], \picorv32_core/n668 );
  and \picorv32_core/sel38_b1/and_b0_2  (\picorv32_core/sel38_b1/B2 , \picorv32_core/latched_rd [1], \picorv32_core/n667 );
  and \picorv32_core/sel38_b1/and_b0_3  (\picorv32_core/sel38_b1/B3 , \picorv32_core/n546 [1], \picorv32_core/n666 );
  and \picorv32_core/sel38_b1/and_b0_4  (\picorv32_core/sel38_b1/B4 , \picorv32_core/latched_rd [1], \picorv32_core/n665 );
  and \picorv32_core/sel38_b1/and_b0_5  (\picorv32_core/sel38_b1/B5 , \picorv32_core/latched_rd [1], \picorv32_core/n664 );
  and \picorv32_core/sel38_b1/and_b0_6  (\picorv32_core/sel38_b1/B6 , \picorv32_core/decoded_rd [1], \picorv32_core/n663 );
  and \picorv32_core/sel38_b1/and_b0_7  (\picorv32_core/sel38_b1/B7 , \picorv32_core/latched_rd [1], \picorv32_core/n662 );
  or \picorv32_core/sel38_b1/or_B0_B1  (\picorv32_core/sel38_b1/or_B0_B1_o , \picorv32_core/sel38_b1/B0 , \picorv32_core/sel38_b1/B1 );
  or \picorv32_core/sel38_b1/or_B2_B3  (\picorv32_core/sel38_b1/or_B2_B3_o , \picorv32_core/sel38_b1/B2 , \picorv32_core/sel38_b1/B3 );
  or \picorv32_core/sel38_b1/or_B4_B5  (\picorv32_core/sel38_b1/or_B4_B5_o , \picorv32_core/sel38_b1/B4 , \picorv32_core/sel38_b1/B5 );
  or \picorv32_core/sel38_b1/or_B6_B7  (\picorv32_core/sel38_b1/or_B6_B7_o , \picorv32_core/sel38_b1/B6 , \picorv32_core/sel38_b1/B7 );
  or \picorv32_core/sel38_b1/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel38_b1/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel38_b1/or_B0_B1_o , \picorv32_core/sel38_b1/or_B2_B3_o );
  or \picorv32_core/sel38_b1/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel38_b1/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel38_b1/or_B4_B5_o , \picorv32_core/sel38_b1/or_B6_B7_o );
  or \picorv32_core/sel38_b1/or_or_or_B0_B1_o_or_  (\picorv32_core/n688 [1], \picorv32_core/sel38_b1/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel38_b1/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel38_b2/and_b0_0  (\picorv32_core/sel38_b2/B0 , \picorv32_core/latched_rd [2], \picorv32_core/n669 );
  and \picorv32_core/sel38_b2/and_b0_1  (\picorv32_core/sel38_b2/B1 , \picorv32_core/latched_rd [2], \picorv32_core/n668 );
  and \picorv32_core/sel38_b2/and_b0_2  (\picorv32_core/sel38_b2/B2 , \picorv32_core/latched_rd [2], \picorv32_core/n667 );
  and \picorv32_core/sel38_b2/and_b0_3  (\picorv32_core/sel38_b2/B3 , \picorv32_core/n546 [2], \picorv32_core/n666 );
  and \picorv32_core/sel38_b2/and_b0_4  (\picorv32_core/sel38_b2/B4 , \picorv32_core/latched_rd [2], \picorv32_core/n665 );
  and \picorv32_core/sel38_b2/and_b0_5  (\picorv32_core/sel38_b2/B5 , \picorv32_core/latched_rd [2], \picorv32_core/n664 );
  and \picorv32_core/sel38_b2/and_b0_6  (\picorv32_core/sel38_b2/B6 , \picorv32_core/decoded_rd [2], \picorv32_core/n663 );
  and \picorv32_core/sel38_b2/and_b0_7  (\picorv32_core/sel38_b2/B7 , \picorv32_core/latched_rd [2], \picorv32_core/n662 );
  or \picorv32_core/sel38_b2/or_B0_B1  (\picorv32_core/sel38_b2/or_B0_B1_o , \picorv32_core/sel38_b2/B0 , \picorv32_core/sel38_b2/B1 );
  or \picorv32_core/sel38_b2/or_B2_B3  (\picorv32_core/sel38_b2/or_B2_B3_o , \picorv32_core/sel38_b2/B2 , \picorv32_core/sel38_b2/B3 );
  or \picorv32_core/sel38_b2/or_B4_B5  (\picorv32_core/sel38_b2/or_B4_B5_o , \picorv32_core/sel38_b2/B4 , \picorv32_core/sel38_b2/B5 );
  or \picorv32_core/sel38_b2/or_B6_B7  (\picorv32_core/sel38_b2/or_B6_B7_o , \picorv32_core/sel38_b2/B6 , \picorv32_core/sel38_b2/B7 );
  or \picorv32_core/sel38_b2/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel38_b2/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel38_b2/or_B0_B1_o , \picorv32_core/sel38_b2/or_B2_B3_o );
  or \picorv32_core/sel38_b2/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel38_b2/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel38_b2/or_B4_B5_o , \picorv32_core/sel38_b2/or_B6_B7_o );
  or \picorv32_core/sel38_b2/or_or_or_B0_B1_o_or_  (\picorv32_core/n688 [2], \picorv32_core/sel38_b2/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel38_b2/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel38_b3/and_b0_0  (\picorv32_core/sel38_b3/B0 , \picorv32_core/latched_rd [3], \picorv32_core/n669 );
  and \picorv32_core/sel38_b3/and_b0_1  (\picorv32_core/sel38_b3/B1 , \picorv32_core/latched_rd [3], \picorv32_core/n668 );
  and \picorv32_core/sel38_b3/and_b0_2  (\picorv32_core/sel38_b3/B2 , \picorv32_core/latched_rd [3], \picorv32_core/n667 );
  and \picorv32_core/sel38_b3/and_b0_3  (\picorv32_core/sel38_b3/B3 , \picorv32_core/n546 [3], \picorv32_core/n666 );
  and \picorv32_core/sel38_b3/and_b0_4  (\picorv32_core/sel38_b3/B4 , \picorv32_core/latched_rd [3], \picorv32_core/n665 );
  and \picorv32_core/sel38_b3/and_b0_5  (\picorv32_core/sel38_b3/B5 , \picorv32_core/latched_rd [3], \picorv32_core/n664 );
  and \picorv32_core/sel38_b3/and_b0_6  (\picorv32_core/sel38_b3/B6 , \picorv32_core/decoded_rd [3], \picorv32_core/n663 );
  and \picorv32_core/sel38_b3/and_b0_7  (\picorv32_core/sel38_b3/B7 , \picorv32_core/latched_rd [3], \picorv32_core/n662 );
  or \picorv32_core/sel38_b3/or_B0_B1  (\picorv32_core/sel38_b3/or_B0_B1_o , \picorv32_core/sel38_b3/B0 , \picorv32_core/sel38_b3/B1 );
  or \picorv32_core/sel38_b3/or_B2_B3  (\picorv32_core/sel38_b3/or_B2_B3_o , \picorv32_core/sel38_b3/B2 , \picorv32_core/sel38_b3/B3 );
  or \picorv32_core/sel38_b3/or_B4_B5  (\picorv32_core/sel38_b3/or_B4_B5_o , \picorv32_core/sel38_b3/B4 , \picorv32_core/sel38_b3/B5 );
  or \picorv32_core/sel38_b3/or_B6_B7  (\picorv32_core/sel38_b3/or_B6_B7_o , \picorv32_core/sel38_b3/B6 , \picorv32_core/sel38_b3/B7 );
  or \picorv32_core/sel38_b3/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel38_b3/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel38_b3/or_B0_B1_o , \picorv32_core/sel38_b3/or_B2_B3_o );
  or \picorv32_core/sel38_b3/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel38_b3/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel38_b3/or_B4_B5_o , \picorv32_core/sel38_b3/or_B6_B7_o );
  or \picorv32_core/sel38_b3/or_or_or_B0_B1_o_or_  (\picorv32_core/n688 [3], \picorv32_core/sel38_b3/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel38_b3/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel38_b4/and_b0_0  (\picorv32_core/sel38_b4/B0 , \picorv32_core/latched_rd [4], \picorv32_core/n669 );
  and \picorv32_core/sel38_b4/and_b0_1  (\picorv32_core/sel38_b4/B1 , \picorv32_core/latched_rd [4], \picorv32_core/n668 );
  and \picorv32_core/sel38_b4/and_b0_2  (\picorv32_core/sel38_b4/B2 , \picorv32_core/latched_rd [4], \picorv32_core/n667 );
  and \picorv32_core/sel38_b4/and_b0_3  (\picorv32_core/sel38_b4/B3 , \picorv32_core/n546 [4], \picorv32_core/n666 );
  and \picorv32_core/sel38_b4/and_b0_4  (\picorv32_core/sel38_b4/B4 , \picorv32_core/latched_rd [4], \picorv32_core/n665 );
  and \picorv32_core/sel38_b4/and_b0_5  (\picorv32_core/sel38_b4/B5 , \picorv32_core/latched_rd [4], \picorv32_core/n664 );
  and \picorv32_core/sel38_b4/and_b0_6  (\picorv32_core/sel38_b4/B6 , \picorv32_core/decoded_rd [4], \picorv32_core/n663 );
  and \picorv32_core/sel38_b4/and_b0_7  (\picorv32_core/sel38_b4/B7 , \picorv32_core/latched_rd [4], \picorv32_core/n662 );
  or \picorv32_core/sel38_b4/or_B0_B1  (\picorv32_core/sel38_b4/or_B0_B1_o , \picorv32_core/sel38_b4/B0 , \picorv32_core/sel38_b4/B1 );
  or \picorv32_core/sel38_b4/or_B2_B3  (\picorv32_core/sel38_b4/or_B2_B3_o , \picorv32_core/sel38_b4/B2 , \picorv32_core/sel38_b4/B3 );
  or \picorv32_core/sel38_b4/or_B4_B5  (\picorv32_core/sel38_b4/or_B4_B5_o , \picorv32_core/sel38_b4/B4 , \picorv32_core/sel38_b4/B5 );
  or \picorv32_core/sel38_b4/or_B6_B7  (\picorv32_core/sel38_b4/or_B6_B7_o , \picorv32_core/sel38_b4/B6 , \picorv32_core/sel38_b4/B7 );
  or \picorv32_core/sel38_b4/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel38_b4/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel38_b4/or_B0_B1_o , \picorv32_core/sel38_b4/or_B2_B3_o );
  or \picorv32_core/sel38_b4/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel38_b4/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel38_b4/or_B4_B5_o , \picorv32_core/sel38_b4/or_B6_B7_o );
  or \picorv32_core/sel38_b4/or_or_or_B0_B1_o_or_  (\picorv32_core/n688 [4], \picorv32_core/sel38_b4/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel38_b4/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel39_b0_sel_is_3  (\picorv32_core/sel39_b0_sel_is_3_o , \picorv32_core/n663 , \picorv32_core/decoder_trigger );
  binary_mux_s3_w1 \picorv32_core/sel3_b0  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [26]),
    .i2(\picorv32_core/mem_rdata_latched [2]),
    .i3(\picorv32_core/n42 [26]),
    .i4(\picorv32_core/n94 [0]),
    .i5(\picorv32_core/n42 [26]),
    .i6(\picorv32_core/mem_rdata_latched [7]),
    .i7(\picorv32_core/n42 [26]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n103 [0]));  // ../src/picorv32.v(504)
  binary_mux_s3_w1 \picorv32_core/sel3_b1  (
    .i0(1'b0),
    .i1(\picorv32_core/n42 [27]),
    .i2(\picorv32_core/mem_rdata_latched [3]),
    .i3(\picorv32_core/n42 [27]),
    .i4(\picorv32_core/n94 [1]),
    .i5(\picorv32_core/n42 [27]),
    .i6(\picorv32_core/mem_rdata_latched [8]),
    .i7(\picorv32_core/n42 [27]),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n103 [1]));  // ../src/picorv32.v(504)
  and \picorv32_core/sel40_b0/and_b0_0  (\picorv32_core/sel40_b0/B0 , \picorv32_core/n661 [0], \picorv32_core/n669 );
  and \picorv32_core/sel40_b0/and_b0_1  (\picorv32_core/sel40_b0/B1 , \picorv32_core/n661 [0], \picorv32_core/n668 );
  and \picorv32_core/sel40_b0/and_b0_2  (\picorv32_core/sel40_b0/B2 , \picorv32_core/n569 [0], \picorv32_core/n667 );
  and \picorv32_core/sel40_b0/and_b0_3  (\picorv32_core/sel40_b0/B3 , \picorv32_core/n549 [0], \picorv32_core/n666 );
  and \picorv32_core/sel40_b0/and_b0_5  (\picorv32_core/sel40_b0/B5 , \picorv32_core/n524 [0], \picorv32_core/n664 );
  and \picorv32_core/sel40_b0/and_b0_6  (\picorv32_core/sel40_b0/B6 , \picorv32_core/n516 [0], \picorv32_core/n663 );
  and \picorv32_core/sel40_b0/and_b0_7  (\picorv32_core/sel40_b0/B7 , \picorv32_core/cpu_state [0], \picorv32_core/n662 );
  or \picorv32_core/sel40_b0/or_B0_B1  (\picorv32_core/sel40_b0/or_B0_B1_o , \picorv32_core/sel40_b0/B0 , \picorv32_core/sel40_b0/B1 );
  or \picorv32_core/sel40_b0/or_B2_B3  (\picorv32_core/sel40_b0/or_B2_B3_o , \picorv32_core/sel40_b0/B2 , \picorv32_core/sel40_b0/B3 );
  or \picorv32_core/sel40_b0/or_B6_B7  (\picorv32_core/sel40_b0/or_B6_B7_o , \picorv32_core/sel40_b0/B6 , \picorv32_core/sel40_b0/B7 );
  or \picorv32_core/sel40_b0/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel40_b0/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b0/or_B0_B1_o , \picorv32_core/sel40_b0/or_B2_B3_o );
  or \picorv32_core/sel40_b0/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel40_b0/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel40_b0/B5 , \picorv32_core/sel40_b0/or_B6_B7_o );
  or \picorv32_core/sel40_b0/or_or_or_B0_B1_o_or_  (\picorv32_core/n692 [0], \picorv32_core/sel40_b0/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b0/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel40_b1/and_b0_0  (\picorv32_core/sel40_b1/B0 , \picorv32_core/n661 [1], \picorv32_core/n669 );
  and \picorv32_core/sel40_b1/and_b0_1  (\picorv32_core/sel40_b1/B1 , \picorv32_core/n661 [1], \picorv32_core/n668 );
  and \picorv32_core/sel40_b1/and_b0_2  (\picorv32_core/sel40_b1/B2 , \picorv32_core/n569 [1], \picorv32_core/n667 );
  and \picorv32_core/sel40_b1/and_b0_3  (\picorv32_core/sel40_b1/B3 , \picorv32_core/n549 [1], \picorv32_core/n666 );
  and \picorv32_core/sel40_b1/and_b0_4  (\picorv32_core/sel40_b1/B4 , \picorv32_core/n521 [1], \picorv32_core/n665 );
  and \picorv32_core/sel40_b1/and_b0_5  (\picorv32_core/sel40_b1/B5 , \picorv32_core/n524 [1], \picorv32_core/n664 );
  and \picorv32_core/sel40_b1/and_b0_6  (\picorv32_core/sel40_b1/B6 , \picorv32_core/n516 [1], \picorv32_core/n663 );
  and \picorv32_core/sel40_b1/and_b0_7  (\picorv32_core/sel40_b1/B7 , \picorv32_core/cpu_state [1], \picorv32_core/n662 );
  or \picorv32_core/sel40_b1/or_B0_B1  (\picorv32_core/sel40_b1/or_B0_B1_o , \picorv32_core/sel40_b1/B0 , \picorv32_core/sel40_b1/B1 );
  or \picorv32_core/sel40_b1/or_B2_B3  (\picorv32_core/sel40_b1/or_B2_B3_o , \picorv32_core/sel40_b1/B2 , \picorv32_core/sel40_b1/B3 );
  or \picorv32_core/sel40_b1/or_B4_B5  (\picorv32_core/sel40_b1/or_B4_B5_o , \picorv32_core/sel40_b1/B4 , \picorv32_core/sel40_b1/B5 );
  or \picorv32_core/sel40_b1/or_B6_B7  (\picorv32_core/sel40_b1/or_B6_B7_o , \picorv32_core/sel40_b1/B6 , \picorv32_core/sel40_b1/B7 );
  or \picorv32_core/sel40_b1/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel40_b1/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b1/or_B0_B1_o , \picorv32_core/sel40_b1/or_B2_B3_o );
  or \picorv32_core/sel40_b1/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel40_b1/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel40_b1/or_B4_B5_o , \picorv32_core/sel40_b1/or_B6_B7_o );
  or \picorv32_core/sel40_b1/or_or_or_B0_B1_o_or_  (\picorv32_core/n692 [1], \picorv32_core/sel40_b1/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b1/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel40_b2/and_b0_0  (\picorv32_core/sel40_b2/B0 , \picorv32_core/n661 [2], \picorv32_core/n669 );
  and \picorv32_core/sel40_b2/and_b0_1  (\picorv32_core/sel40_b2/B1 , \picorv32_core/n661 [2], \picorv32_core/n668 );
  and \picorv32_core/sel40_b2/and_b0_2  (\picorv32_core/sel40_b2/B2 , \picorv32_core/n569 [2], \picorv32_core/n667 );
  and \picorv32_core/sel40_b2/and_b0_3  (\picorv32_core/sel40_b2/B3 , \picorv32_core/n549 [2], \picorv32_core/n666 );
  and \picorv32_core/sel40_b2/and_b0_4  (\picorv32_core/sel40_b2/B4 , \picorv32_core/n521 [2], \picorv32_core/n665 );
  and \picorv32_core/sel40_b2/and_b0_5  (\picorv32_core/sel40_b2/B5 , \picorv32_core/sel19_b2/or_B0_or_B1_B2_o_o , \picorv32_core/n664 );
  and \picorv32_core/sel40_b2/and_b0_6  (\picorv32_core/sel40_b2/B6 , \picorv32_core/n516 [2], \picorv32_core/n663 );
  and \picorv32_core/sel40_b2/and_b0_7  (\picorv32_core/sel40_b2/B7 , \picorv32_core/cpu_state [2], \picorv32_core/n662 );
  or \picorv32_core/sel40_b2/or_B0_B1  (\picorv32_core/sel40_b2/or_B0_B1_o , \picorv32_core/sel40_b2/B0 , \picorv32_core/sel40_b2/B1 );
  or \picorv32_core/sel40_b2/or_B2_B3  (\picorv32_core/sel40_b2/or_B2_B3_o , \picorv32_core/sel40_b2/B2 , \picorv32_core/sel40_b2/B3 );
  or \picorv32_core/sel40_b2/or_B4_B5  (\picorv32_core/sel40_b2/or_B4_B5_o , \picorv32_core/sel40_b2/B4 , \picorv32_core/sel40_b2/B5 );
  or \picorv32_core/sel40_b2/or_B6_B7  (\picorv32_core/sel40_b2/or_B6_B7_o , \picorv32_core/sel40_b2/B6 , \picorv32_core/sel40_b2/B7 );
  or \picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b2/or_B0_B1_o , \picorv32_core/sel40_b2/or_B2_B3_o );
  or \picorv32_core/sel40_b2/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel40_b2/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel40_b2/or_B4_B5_o , \picorv32_core/sel40_b2/or_B6_B7_o );
  or \picorv32_core/sel40_b2/or_or_or_B0_B1_o_or_  (\picorv32_core/n692 [2], \picorv32_core/sel40_b2/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b2/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel40_b3/and_b0_0  (\picorv32_core/sel40_b3/B0 , \picorv32_core/n661 [3], \picorv32_core/n669 );
  and \picorv32_core/sel40_b3/and_b0_1  (\picorv32_core/sel40_b3/B1 , \picorv32_core/n661 [3], \picorv32_core/n668 );
  and \picorv32_core/sel40_b3/and_b0_2  (\picorv32_core/sel40_b3/B2 , \picorv32_core/n569 [3], \picorv32_core/n667 );
  and \picorv32_core/sel40_b3/and_b0_3  (\picorv32_core/sel40_b3/B3 , \picorv32_core/n549 [3], \picorv32_core/n666 );
  and \picorv32_core/sel40_b3/and_b0_4  (\picorv32_core/sel40_b3/B4 , \picorv32_core/n521 [3], \picorv32_core/n665 );
  and \picorv32_core/sel40_b3/and_b0_5  (\picorv32_core/sel40_b3/B5 , \picorv32_core/n524 [3], \picorv32_core/n664 );
  and \picorv32_core/sel40_b3/and_b0_6  (\picorv32_core/sel40_b3/B6 , \picorv32_core/n516 [3], \picorv32_core/n663 );
  and \picorv32_core/sel40_b3/and_b0_7  (\picorv32_core/sel40_b3/B7 , \picorv32_core/cpu_state [3], \picorv32_core/n662 );
  or \picorv32_core/sel40_b3/or_B0_B1  (\picorv32_core/sel40_b3/or_B0_B1_o , \picorv32_core/sel40_b3/B0 , \picorv32_core/sel40_b3/B1 );
  or \picorv32_core/sel40_b3/or_B2_B3  (\picorv32_core/sel40_b3/or_B2_B3_o , \picorv32_core/sel40_b3/B2 , \picorv32_core/sel40_b3/B3 );
  or \picorv32_core/sel40_b3/or_B4_B5  (\picorv32_core/sel40_b3/or_B4_B5_o , \picorv32_core/sel40_b3/B4 , \picorv32_core/sel40_b3/B5 );
  or \picorv32_core/sel40_b3/or_B6_B7  (\picorv32_core/sel40_b3/or_B6_B7_o , \picorv32_core/sel40_b3/B6 , \picorv32_core/sel40_b3/B7 );
  or \picorv32_core/sel40_b3/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel40_b3/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b3/or_B0_B1_o , \picorv32_core/sel40_b3/or_B2_B3_o );
  or \picorv32_core/sel40_b3/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel40_b3/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel40_b3/or_B4_B5_o , \picorv32_core/sel40_b3/or_B6_B7_o );
  or \picorv32_core/sel40_b3/or_or_or_B0_B1_o_or_  (\picorv32_core/n692 [3], \picorv32_core/sel40_b3/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b3/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel40_b4/and_b0_0  (\picorv32_core/sel40_b4/B0 , \picorv32_core/n661 [4], \picorv32_core/n669 );
  and \picorv32_core/sel40_b4/and_b0_1  (\picorv32_core/sel40_b4/B1 , \picorv32_core/n661 [4], \picorv32_core/n668 );
  and \picorv32_core/sel40_b4/and_b0_2  (\picorv32_core/sel40_b4/B2 , \picorv32_core/n569 [4], \picorv32_core/n667 );
  and \picorv32_core/sel40_b4/and_b0_3  (\picorv32_core/sel40_b4/B3 , \picorv32_core/n549 [4], \picorv32_core/n666 );
  and \picorv32_core/sel40_b4/and_b0_6  (\picorv32_core/sel40_b4/B6 , \picorv32_core/n516 [4], \picorv32_core/n663 );
  and \picorv32_core/sel40_b4/and_b0_7  (\picorv32_core/sel40_b4/B7 , \picorv32_core/cpu_state [4], \picorv32_core/n662 );
  or \picorv32_core/sel40_b4/or_B0_B1  (\picorv32_core/sel40_b4/or_B0_B1_o , \picorv32_core/sel40_b4/B0 , \picorv32_core/sel40_b4/B1 );
  or \picorv32_core/sel40_b4/or_B2_B3  (\picorv32_core/sel40_b4/or_B2_B3_o , \picorv32_core/sel40_b4/B2 , \picorv32_core/sel40_b4/B3 );
  or \picorv32_core/sel40_b4/or_B6_B7  (\picorv32_core/sel40_b4/or_B6_B7_o , \picorv32_core/sel40_b4/B6 , \picorv32_core/sel40_b4/B7 );
  or \picorv32_core/sel40_b4/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel40_b4/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b4/or_B0_B1_o , \picorv32_core/sel40_b4/or_B2_B3_o );
  or \picorv32_core/sel40_b4/or_or_or_B0_B1_o_or_  (\picorv32_core/n692 [4], \picorv32_core/sel40_b4/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b4/or_B6_B7_o );
  and \picorv32_core/sel40_b5/and_b0_0  (\picorv32_core/sel40_b5/B0 , \picorv32_core/n661 [5], \picorv32_core/n669 );
  and \picorv32_core/sel40_b5/and_b0_1  (\picorv32_core/sel40_b5/B1 , \picorv32_core/n661 [5], \picorv32_core/n668 );
  and \picorv32_core/sel40_b5/and_b0_2  (\picorv32_core/sel40_b5/B2 , \picorv32_core/n569 [5], \picorv32_core/n667 );
  and \picorv32_core/sel40_b5/and_b0_3  (\picorv32_core/sel40_b5/B3 , \picorv32_core/n549 [5], \picorv32_core/n666 );
  and \picorv32_core/sel40_b5/and_b0_6  (\picorv32_core/sel40_b5/B6 , \picorv32_core/n516 [5], \picorv32_core/n663 );
  and \picorv32_core/sel40_b5/and_b0_7  (\picorv32_core/sel40_b5/B7 , \picorv32_core/cpu_state [5], \picorv32_core/n662 );
  or \picorv32_core/sel40_b5/or_B0_B1  (\picorv32_core/sel40_b5/or_B0_B1_o , \picorv32_core/sel40_b5/B0 , \picorv32_core/sel40_b5/B1 );
  or \picorv32_core/sel40_b5/or_B2_B3  (\picorv32_core/sel40_b5/or_B2_B3_o , \picorv32_core/sel40_b5/B2 , \picorv32_core/sel40_b5/B3 );
  or \picorv32_core/sel40_b5/or_B6_B7  (\picorv32_core/sel40_b5/or_B6_B7_o , \picorv32_core/sel40_b5/B6 , \picorv32_core/sel40_b5/B7 );
  or \picorv32_core/sel40_b5/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel40_b5/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b5/or_B0_B1_o , \picorv32_core/sel40_b5/or_B2_B3_o );
  or \picorv32_core/sel40_b5/or_or_or_B0_B1_o_or_  (\picorv32_core/n692 [5], \picorv32_core/sel40_b5/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b5/or_B6_B7_o );
  and \picorv32_core/sel40_b6/and_b0_0  (\picorv32_core/sel40_b6/B0 , \picorv32_core/n661 [6], \picorv32_core/n669 );
  and \picorv32_core/sel40_b6/and_b0_1  (\picorv32_core/sel40_b6/B1 , \picorv32_core/n661 [6], \picorv32_core/n668 );
  and \picorv32_core/sel40_b6/and_b0_2  (\picorv32_core/sel40_b6/B2 , \picorv32_core/n569 [6], \picorv32_core/n667 );
  and \picorv32_core/sel40_b6/and_b0_3  (\picorv32_core/sel40_b6/B3 , \picorv32_core/n549 [6], \picorv32_core/n666 );
  and \picorv32_core/sel40_b6/and_b0_5  (\picorv32_core/sel40_b6/B5 , \picorv32_core/n524 [6], \picorv32_core/n664 );
  and \picorv32_core/sel40_b6/and_b0_6  (\picorv32_core/sel40_b6/B6 , \picorv32_core/n516 [6], \picorv32_core/n663 );
  and \picorv32_core/sel40_b6/and_b0_7  (\picorv32_core/sel40_b6/B7 , \picorv32_core/cpu_state [6], \picorv32_core/n662 );
  or \picorv32_core/sel40_b6/or_B0_B1  (\picorv32_core/sel40_b6/or_B0_B1_o , \picorv32_core/sel40_b6/B0 , \picorv32_core/sel40_b6/B1 );
  or \picorv32_core/sel40_b6/or_B2_B3  (\picorv32_core/sel40_b6/or_B2_B3_o , \picorv32_core/sel40_b6/B2 , \picorv32_core/sel40_b6/B3 );
  or \picorv32_core/sel40_b6/or_B6_B7  (\picorv32_core/sel40_b6/or_B6_B7_o , \picorv32_core/sel40_b6/B6 , \picorv32_core/sel40_b6/B7 );
  or \picorv32_core/sel40_b6/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel40_b6/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b6/or_B0_B1_o , \picorv32_core/sel40_b6/or_B2_B3_o );
  or \picorv32_core/sel40_b6/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel40_b6/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel40_b6/B5 , \picorv32_core/sel40_b6/or_B6_B7_o );
  or \picorv32_core/sel40_b6/or_or_or_B0_B1_o_or_  (\picorv32_core/n692 [6], \picorv32_core/sel40_b6/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b6/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel40_b7/and_b0_0  (\picorv32_core/sel40_b7/B0 , \picorv32_core/n661 [7], \picorv32_core/n669 );
  and \picorv32_core/sel40_b7/and_b0_1  (\picorv32_core/sel40_b7/B1 , \picorv32_core/n661 [7], \picorv32_core/n668 );
  and \picorv32_core/sel40_b7/and_b0_2  (\picorv32_core/sel40_b7/B2 , \picorv32_core/n569 [7], \picorv32_core/n667 );
  and \picorv32_core/sel40_b7/and_b0_3  (\picorv32_core/sel40_b7/B3 , \picorv32_core/n549 [7], \picorv32_core/n666 );
  and \picorv32_core/sel40_b7/and_b0_5  (\picorv32_core/sel40_b7/B5 , \picorv32_core/n524 [7], \picorv32_core/n664 );
  and \picorv32_core/sel40_b7/and_b0_6  (\picorv32_core/sel40_b7/B6 , \picorv32_core/n516 [7], \picorv32_core/n663 );
  and \picorv32_core/sel40_b7/and_b0_7  (\picorv32_core/sel40_b7/B7 , \picorv32_core/cpu_state [7], \picorv32_core/n662 );
  or \picorv32_core/sel40_b7/or_B0_B1  (\picorv32_core/sel40_b7/or_B0_B1_o , \picorv32_core/sel40_b7/B0 , \picorv32_core/sel40_b7/B1 );
  or \picorv32_core/sel40_b7/or_B2_B3  (\picorv32_core/sel40_b7/or_B2_B3_o , \picorv32_core/sel40_b7/B2 , \picorv32_core/sel40_b7/B3 );
  or \picorv32_core/sel40_b7/or_B6_B7  (\picorv32_core/sel40_b7/or_B6_B7_o , \picorv32_core/sel40_b7/B6 , \picorv32_core/sel40_b7/B7 );
  or \picorv32_core/sel40_b7/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel40_b7/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b7/or_B0_B1_o , \picorv32_core/sel40_b7/or_B2_B3_o );
  or \picorv32_core/sel40_b7/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel40_b7/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel40_b7/B5 , \picorv32_core/sel40_b7/or_B6_B7_o );
  or \picorv32_core/sel40_b7/or_or_or_B0_B1_o_or_  (\picorv32_core/n692 [7], \picorv32_core/sel40_b7/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel40_b7/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b0/and_b0_0  (\picorv32_core/sel41_b0/B0 , \picorv32_core/n656 [0], \picorv32_core/n669 );
  and \picorv32_core/sel41_b0/and_b0_1  (\picorv32_core/sel41_b0/B1 , \picorv32_core/n584 [0], \picorv32_core/n668 );
  and \picorv32_core/sel41_b0/and_b0_2  (\picorv32_core/sel41_b0/B2 , \picorv32_core/n570 [0], \picorv32_core/n667 );
  and \picorv32_core/sel41_b0/and_b0_3  (\picorv32_core/sel41_b0/B3 , \picorv32_core/pcpi_rs1$0$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b0/and_b0_4  (\picorv32_core/sel41_b0/B4 , \picorv32_core/pcpi_rs1$0$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b0/and_b0_5  (\picorv32_core/sel41_b0/B5 , \picorv32_core/n527 [0], \picorv32_core/n664 );
  and \picorv32_core/sel41_b0/and_b0_6  (\picorv32_core/sel41_b0/B6 , \picorv32_core/pcpi_rs1$0$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b0/and_b0_7  (\picorv32_core/sel41_b0/B7 , \picorv32_core/pcpi_rs1$0$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b0/or_B0_B1  (\picorv32_core/sel41_b0/or_B0_B1_o , \picorv32_core/sel41_b0/B0 , \picorv32_core/sel41_b0/B1 );
  or \picorv32_core/sel41_b0/or_B2_B3  (\picorv32_core/sel41_b0/or_B2_B3_o , \picorv32_core/sel41_b0/B2 , \picorv32_core/sel41_b0/B3 );
  or \picorv32_core/sel41_b0/or_B4_B5  (\picorv32_core/sel41_b0/or_B4_B5_o , \picorv32_core/sel41_b0/B4 , \picorv32_core/sel41_b0/B5 );
  or \picorv32_core/sel41_b0/or_B6_B7  (\picorv32_core/sel41_b0/or_B6_B7_o , \picorv32_core/sel41_b0/B6 , \picorv32_core/sel41_b0/B7 );
  or \picorv32_core/sel41_b0/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b0/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b0/or_B0_B1_o , \picorv32_core/sel41_b0/or_B2_B3_o );
  or \picorv32_core/sel41_b0/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b0/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b0/or_B4_B5_o , \picorv32_core/sel41_b0/or_B6_B7_o );
  or \picorv32_core/sel41_b0/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [0], \picorv32_core/sel41_b0/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b0/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b1/and_b0_0  (\picorv32_core/sel41_b1/B0 , \picorv32_core/n656 [1], \picorv32_core/n669 );
  and \picorv32_core/sel41_b1/and_b0_1  (\picorv32_core/sel41_b1/B1 , \picorv32_core/n584 [1], \picorv32_core/n668 );
  and \picorv32_core/sel41_b1/and_b0_2  (\picorv32_core/sel41_b1/B2 , \picorv32_core/n570 [1], \picorv32_core/n667 );
  and \picorv32_core/sel41_b1/and_b0_3  (\picorv32_core/sel41_b1/B3 , \picorv32_core/pcpi_rs1$1$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b1/and_b0_4  (\picorv32_core/sel41_b1/B4 , \picorv32_core/pcpi_rs1$1$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b1/and_b0_5  (\picorv32_core/sel41_b1/B5 , \picorv32_core/n527 [1], \picorv32_core/n664 );
  and \picorv32_core/sel41_b1/and_b0_6  (\picorv32_core/sel41_b1/B6 , \picorv32_core/pcpi_rs1$1$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b1/and_b0_7  (\picorv32_core/sel41_b1/B7 , \picorv32_core/pcpi_rs1$1$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b1/or_B0_B1  (\picorv32_core/sel41_b1/or_B0_B1_o , \picorv32_core/sel41_b1/B0 , \picorv32_core/sel41_b1/B1 );
  or \picorv32_core/sel41_b1/or_B2_B3  (\picorv32_core/sel41_b1/or_B2_B3_o , \picorv32_core/sel41_b1/B2 , \picorv32_core/sel41_b1/B3 );
  or \picorv32_core/sel41_b1/or_B4_B5  (\picorv32_core/sel41_b1/or_B4_B5_o , \picorv32_core/sel41_b1/B4 , \picorv32_core/sel41_b1/B5 );
  or \picorv32_core/sel41_b1/or_B6_B7  (\picorv32_core/sel41_b1/or_B6_B7_o , \picorv32_core/sel41_b1/B6 , \picorv32_core/sel41_b1/B7 );
  or \picorv32_core/sel41_b1/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b1/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b1/or_B0_B1_o , \picorv32_core/sel41_b1/or_B2_B3_o );
  or \picorv32_core/sel41_b1/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b1/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b1/or_B4_B5_o , \picorv32_core/sel41_b1/or_B6_B7_o );
  or \picorv32_core/sel41_b1/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [1], \picorv32_core/sel41_b1/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b1/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b10/and_b0_0  (\picorv32_core/sel41_b10/B0 , \picorv32_core/n656 [10], \picorv32_core/n669 );
  and \picorv32_core/sel41_b10/and_b0_1  (\picorv32_core/sel41_b10/B1 , \picorv32_core/n584 [10], \picorv32_core/n668 );
  and \picorv32_core/sel41_b10/and_b0_2  (\picorv32_core/sel41_b10/B2 , \picorv32_core/n570 [10], \picorv32_core/n667 );
  and \picorv32_core/sel41_b10/and_b0_3  (\picorv32_core/sel41_b10/B3 , \picorv32_core/pcpi_rs1$10$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b10/and_b0_4  (\picorv32_core/sel41_b10/B4 , \picorv32_core/pcpi_rs1$10$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b10/and_b0_5  (\picorv32_core/sel41_b10/B5 , \picorv32_core/n527 [10], \picorv32_core/n664 );
  and \picorv32_core/sel41_b10/and_b0_6  (\picorv32_core/sel41_b10/B6 , \picorv32_core/pcpi_rs1$10$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b10/and_b0_7  (\picorv32_core/sel41_b10/B7 , \picorv32_core/pcpi_rs1$10$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b10/or_B0_B1  (\picorv32_core/sel41_b10/or_B0_B1_o , \picorv32_core/sel41_b10/B0 , \picorv32_core/sel41_b10/B1 );
  or \picorv32_core/sel41_b10/or_B2_B3  (\picorv32_core/sel41_b10/or_B2_B3_o , \picorv32_core/sel41_b10/B2 , \picorv32_core/sel41_b10/B3 );
  or \picorv32_core/sel41_b10/or_B4_B5  (\picorv32_core/sel41_b10/or_B4_B5_o , \picorv32_core/sel41_b10/B4 , \picorv32_core/sel41_b10/B5 );
  or \picorv32_core/sel41_b10/or_B6_B7  (\picorv32_core/sel41_b10/or_B6_B7_o , \picorv32_core/sel41_b10/B6 , \picorv32_core/sel41_b10/B7 );
  or \picorv32_core/sel41_b10/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b10/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b10/or_B0_B1_o , \picorv32_core/sel41_b10/or_B2_B3_o );
  or \picorv32_core/sel41_b10/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b10/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b10/or_B4_B5_o , \picorv32_core/sel41_b10/or_B6_B7_o );
  or \picorv32_core/sel41_b10/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [10], \picorv32_core/sel41_b10/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b10/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b11/and_b0_0  (\picorv32_core/sel41_b11/B0 , \picorv32_core/n656 [11], \picorv32_core/n669 );
  and \picorv32_core/sel41_b11/and_b0_1  (\picorv32_core/sel41_b11/B1 , \picorv32_core/n584 [11], \picorv32_core/n668 );
  and \picorv32_core/sel41_b11/and_b0_2  (\picorv32_core/sel41_b11/B2 , \picorv32_core/n570 [11], \picorv32_core/n667 );
  and \picorv32_core/sel41_b11/and_b0_3  (\picorv32_core/sel41_b11/B3 , \picorv32_core/pcpi_rs1$11$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b11/and_b0_4  (\picorv32_core/sel41_b11/B4 , \picorv32_core/pcpi_rs1$11$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b11/and_b0_5  (\picorv32_core/sel41_b11/B5 , \picorv32_core/n527 [11], \picorv32_core/n664 );
  and \picorv32_core/sel41_b11/and_b0_6  (\picorv32_core/sel41_b11/B6 , \picorv32_core/pcpi_rs1$11$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b11/and_b0_7  (\picorv32_core/sel41_b11/B7 , \picorv32_core/pcpi_rs1$11$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b11/or_B0_B1  (\picorv32_core/sel41_b11/or_B0_B1_o , \picorv32_core/sel41_b11/B0 , \picorv32_core/sel41_b11/B1 );
  or \picorv32_core/sel41_b11/or_B2_B3  (\picorv32_core/sel41_b11/or_B2_B3_o , \picorv32_core/sel41_b11/B2 , \picorv32_core/sel41_b11/B3 );
  or \picorv32_core/sel41_b11/or_B4_B5  (\picorv32_core/sel41_b11/or_B4_B5_o , \picorv32_core/sel41_b11/B4 , \picorv32_core/sel41_b11/B5 );
  or \picorv32_core/sel41_b11/or_B6_B7  (\picorv32_core/sel41_b11/or_B6_B7_o , \picorv32_core/sel41_b11/B6 , \picorv32_core/sel41_b11/B7 );
  or \picorv32_core/sel41_b11/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b11/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b11/or_B0_B1_o , \picorv32_core/sel41_b11/or_B2_B3_o );
  or \picorv32_core/sel41_b11/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b11/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b11/or_B4_B5_o , \picorv32_core/sel41_b11/or_B6_B7_o );
  or \picorv32_core/sel41_b11/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [11], \picorv32_core/sel41_b11/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b11/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b12/and_b0_0  (\picorv32_core/sel41_b12/B0 , \picorv32_core/n656 [12], \picorv32_core/n669 );
  and \picorv32_core/sel41_b12/and_b0_1  (\picorv32_core/sel41_b12/B1 , \picorv32_core/n584 [12], \picorv32_core/n668 );
  and \picorv32_core/sel41_b12/and_b0_2  (\picorv32_core/sel41_b12/B2 , \picorv32_core/n570 [12], \picorv32_core/n667 );
  and \picorv32_core/sel41_b12/and_b0_3  (\picorv32_core/sel41_b12/B3 , \picorv32_core/pcpi_rs1$12$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b12/and_b0_4  (\picorv32_core/sel41_b12/B4 , \picorv32_core/pcpi_rs1$12$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b12/and_b0_5  (\picorv32_core/sel41_b12/B5 , \picorv32_core/n527 [12], \picorv32_core/n664 );
  and \picorv32_core/sel41_b12/and_b0_6  (\picorv32_core/sel41_b12/B6 , \picorv32_core/pcpi_rs1$12$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b12/and_b0_7  (\picorv32_core/sel41_b12/B7 , \picorv32_core/pcpi_rs1$12$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b12/or_B0_B1  (\picorv32_core/sel41_b12/or_B0_B1_o , \picorv32_core/sel41_b12/B0 , \picorv32_core/sel41_b12/B1 );
  or \picorv32_core/sel41_b12/or_B2_B3  (\picorv32_core/sel41_b12/or_B2_B3_o , \picorv32_core/sel41_b12/B2 , \picorv32_core/sel41_b12/B3 );
  or \picorv32_core/sel41_b12/or_B4_B5  (\picorv32_core/sel41_b12/or_B4_B5_o , \picorv32_core/sel41_b12/B4 , \picorv32_core/sel41_b12/B5 );
  or \picorv32_core/sel41_b12/or_B6_B7  (\picorv32_core/sel41_b12/or_B6_B7_o , \picorv32_core/sel41_b12/B6 , \picorv32_core/sel41_b12/B7 );
  or \picorv32_core/sel41_b12/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b12/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b12/or_B0_B1_o , \picorv32_core/sel41_b12/or_B2_B3_o );
  or \picorv32_core/sel41_b12/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b12/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b12/or_B4_B5_o , \picorv32_core/sel41_b12/or_B6_B7_o );
  or \picorv32_core/sel41_b12/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [12], \picorv32_core/sel41_b12/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b12/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b13/and_b0_0  (\picorv32_core/sel41_b13/B0 , \picorv32_core/n656 [13], \picorv32_core/n669 );
  and \picorv32_core/sel41_b13/and_b0_1  (\picorv32_core/sel41_b13/B1 , \picorv32_core/n584 [13], \picorv32_core/n668 );
  and \picorv32_core/sel41_b13/and_b0_2  (\picorv32_core/sel41_b13/B2 , \picorv32_core/n570 [13], \picorv32_core/n667 );
  and \picorv32_core/sel41_b13/and_b0_3  (\picorv32_core/sel41_b13/B3 , \picorv32_core/pcpi_rs1$13$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b13/and_b0_4  (\picorv32_core/sel41_b13/B4 , \picorv32_core/pcpi_rs1$13$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b13/and_b0_5  (\picorv32_core/sel41_b13/B5 , \picorv32_core/n527 [13], \picorv32_core/n664 );
  and \picorv32_core/sel41_b13/and_b0_6  (\picorv32_core/sel41_b13/B6 , \picorv32_core/pcpi_rs1$13$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b13/and_b0_7  (\picorv32_core/sel41_b13/B7 , \picorv32_core/pcpi_rs1$13$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b13/or_B0_B1  (\picorv32_core/sel41_b13/or_B0_B1_o , \picorv32_core/sel41_b13/B0 , \picorv32_core/sel41_b13/B1 );
  or \picorv32_core/sel41_b13/or_B2_B3  (\picorv32_core/sel41_b13/or_B2_B3_o , \picorv32_core/sel41_b13/B2 , \picorv32_core/sel41_b13/B3 );
  or \picorv32_core/sel41_b13/or_B4_B5  (\picorv32_core/sel41_b13/or_B4_B5_o , \picorv32_core/sel41_b13/B4 , \picorv32_core/sel41_b13/B5 );
  or \picorv32_core/sel41_b13/or_B6_B7  (\picorv32_core/sel41_b13/or_B6_B7_o , \picorv32_core/sel41_b13/B6 , \picorv32_core/sel41_b13/B7 );
  or \picorv32_core/sel41_b13/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b13/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b13/or_B0_B1_o , \picorv32_core/sel41_b13/or_B2_B3_o );
  or \picorv32_core/sel41_b13/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b13/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b13/or_B4_B5_o , \picorv32_core/sel41_b13/or_B6_B7_o );
  or \picorv32_core/sel41_b13/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [13], \picorv32_core/sel41_b13/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b13/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b14/and_b0_0  (\picorv32_core/sel41_b14/B0 , \picorv32_core/n656 [14], \picorv32_core/n669 );
  and \picorv32_core/sel41_b14/and_b0_1  (\picorv32_core/sel41_b14/B1 , \picorv32_core/n584 [14], \picorv32_core/n668 );
  and \picorv32_core/sel41_b14/and_b0_2  (\picorv32_core/sel41_b14/B2 , \picorv32_core/n570 [14], \picorv32_core/n667 );
  and \picorv32_core/sel41_b14/and_b0_3  (\picorv32_core/sel41_b14/B3 , \picorv32_core/pcpi_rs1$14$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b14/and_b0_4  (\picorv32_core/sel41_b14/B4 , \picorv32_core/pcpi_rs1$14$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b14/and_b0_5  (\picorv32_core/sel41_b14/B5 , \picorv32_core/n527 [14], \picorv32_core/n664 );
  and \picorv32_core/sel41_b14/and_b0_6  (\picorv32_core/sel41_b14/B6 , \picorv32_core/pcpi_rs1$14$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b14/and_b0_7  (\picorv32_core/sel41_b14/B7 , \picorv32_core/pcpi_rs1$14$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b14/or_B0_B1  (\picorv32_core/sel41_b14/or_B0_B1_o , \picorv32_core/sel41_b14/B0 , \picorv32_core/sel41_b14/B1 );
  or \picorv32_core/sel41_b14/or_B2_B3  (\picorv32_core/sel41_b14/or_B2_B3_o , \picorv32_core/sel41_b14/B2 , \picorv32_core/sel41_b14/B3 );
  or \picorv32_core/sel41_b14/or_B4_B5  (\picorv32_core/sel41_b14/or_B4_B5_o , \picorv32_core/sel41_b14/B4 , \picorv32_core/sel41_b14/B5 );
  or \picorv32_core/sel41_b14/or_B6_B7  (\picorv32_core/sel41_b14/or_B6_B7_o , \picorv32_core/sel41_b14/B6 , \picorv32_core/sel41_b14/B7 );
  or \picorv32_core/sel41_b14/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b14/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b14/or_B0_B1_o , \picorv32_core/sel41_b14/or_B2_B3_o );
  or \picorv32_core/sel41_b14/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b14/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b14/or_B4_B5_o , \picorv32_core/sel41_b14/or_B6_B7_o );
  or \picorv32_core/sel41_b14/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [14], \picorv32_core/sel41_b14/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b14/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b15/and_b0_0  (\picorv32_core/sel41_b15/B0 , \picorv32_core/n656 [15], \picorv32_core/n669 );
  and \picorv32_core/sel41_b15/and_b0_1  (\picorv32_core/sel41_b15/B1 , \picorv32_core/n584 [15], \picorv32_core/n668 );
  and \picorv32_core/sel41_b15/and_b0_2  (\picorv32_core/sel41_b15/B2 , \picorv32_core/n570 [15], \picorv32_core/n667 );
  and \picorv32_core/sel41_b15/and_b0_3  (\picorv32_core/sel41_b15/B3 , \picorv32_core/pcpi_rs1$15$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b15/and_b0_4  (\picorv32_core/sel41_b15/B4 , \picorv32_core/pcpi_rs1$15$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b15/and_b0_5  (\picorv32_core/sel41_b15/B5 , \picorv32_core/n527 [15], \picorv32_core/n664 );
  and \picorv32_core/sel41_b15/and_b0_6  (\picorv32_core/sel41_b15/B6 , \picorv32_core/pcpi_rs1$15$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b15/and_b0_7  (\picorv32_core/sel41_b15/B7 , \picorv32_core/pcpi_rs1$15$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b15/or_B0_B1  (\picorv32_core/sel41_b15/or_B0_B1_o , \picorv32_core/sel41_b15/B0 , \picorv32_core/sel41_b15/B1 );
  or \picorv32_core/sel41_b15/or_B2_B3  (\picorv32_core/sel41_b15/or_B2_B3_o , \picorv32_core/sel41_b15/B2 , \picorv32_core/sel41_b15/B3 );
  or \picorv32_core/sel41_b15/or_B4_B5  (\picorv32_core/sel41_b15/or_B4_B5_o , \picorv32_core/sel41_b15/B4 , \picorv32_core/sel41_b15/B5 );
  or \picorv32_core/sel41_b15/or_B6_B7  (\picorv32_core/sel41_b15/or_B6_B7_o , \picorv32_core/sel41_b15/B6 , \picorv32_core/sel41_b15/B7 );
  or \picorv32_core/sel41_b15/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b15/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b15/or_B0_B1_o , \picorv32_core/sel41_b15/or_B2_B3_o );
  or \picorv32_core/sel41_b15/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b15/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b15/or_B4_B5_o , \picorv32_core/sel41_b15/or_B6_B7_o );
  or \picorv32_core/sel41_b15/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [15], \picorv32_core/sel41_b15/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b15/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b16/and_b0_0  (\picorv32_core/sel41_b16/B0 , \picorv32_core/n656 [16], \picorv32_core/n669 );
  and \picorv32_core/sel41_b16/and_b0_1  (\picorv32_core/sel41_b16/B1 , \picorv32_core/n584 [16], \picorv32_core/n668 );
  and \picorv32_core/sel41_b16/and_b0_2  (\picorv32_core/sel41_b16/B2 , \picorv32_core/n570 [16], \picorv32_core/n667 );
  and \picorv32_core/sel41_b16/and_b0_3  (\picorv32_core/sel41_b16/B3 , \picorv32_core/pcpi_rs1$16$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b16/and_b0_4  (\picorv32_core/sel41_b16/B4 , \picorv32_core/pcpi_rs1$16$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b16/and_b0_5  (\picorv32_core/sel41_b16/B5 , \picorv32_core/n527 [16], \picorv32_core/n664 );
  and \picorv32_core/sel41_b16/and_b0_6  (\picorv32_core/sel41_b16/B6 , \picorv32_core/pcpi_rs1$16$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b16/and_b0_7  (\picorv32_core/sel41_b16/B7 , \picorv32_core/pcpi_rs1$16$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b16/or_B0_B1  (\picorv32_core/sel41_b16/or_B0_B1_o , \picorv32_core/sel41_b16/B0 , \picorv32_core/sel41_b16/B1 );
  or \picorv32_core/sel41_b16/or_B2_B3  (\picorv32_core/sel41_b16/or_B2_B3_o , \picorv32_core/sel41_b16/B2 , \picorv32_core/sel41_b16/B3 );
  or \picorv32_core/sel41_b16/or_B4_B5  (\picorv32_core/sel41_b16/or_B4_B5_o , \picorv32_core/sel41_b16/B4 , \picorv32_core/sel41_b16/B5 );
  or \picorv32_core/sel41_b16/or_B6_B7  (\picorv32_core/sel41_b16/or_B6_B7_o , \picorv32_core/sel41_b16/B6 , \picorv32_core/sel41_b16/B7 );
  or \picorv32_core/sel41_b16/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b16/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b16/or_B0_B1_o , \picorv32_core/sel41_b16/or_B2_B3_o );
  or \picorv32_core/sel41_b16/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b16/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b16/or_B4_B5_o , \picorv32_core/sel41_b16/or_B6_B7_o );
  or \picorv32_core/sel41_b16/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [16], \picorv32_core/sel41_b16/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b16/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b17/and_b0_0  (\picorv32_core/sel41_b17/B0 , \picorv32_core/n656 [17], \picorv32_core/n669 );
  and \picorv32_core/sel41_b17/and_b0_1  (\picorv32_core/sel41_b17/B1 , \picorv32_core/n584 [17], \picorv32_core/n668 );
  and \picorv32_core/sel41_b17/and_b0_2  (\picorv32_core/sel41_b17/B2 , \picorv32_core/n570 [17], \picorv32_core/n667 );
  and \picorv32_core/sel41_b17/and_b0_3  (\picorv32_core/sel41_b17/B3 , \picorv32_core/pcpi_rs1$17$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b17/and_b0_4  (\picorv32_core/sel41_b17/B4 , \picorv32_core/pcpi_rs1$17$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b17/and_b0_5  (\picorv32_core/sel41_b17/B5 , \picorv32_core/n527 [17], \picorv32_core/n664 );
  and \picorv32_core/sel41_b17/and_b0_6  (\picorv32_core/sel41_b17/B6 , \picorv32_core/pcpi_rs1$17$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b17/and_b0_7  (\picorv32_core/sel41_b17/B7 , \picorv32_core/pcpi_rs1$17$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b17/or_B0_B1  (\picorv32_core/sel41_b17/or_B0_B1_o , \picorv32_core/sel41_b17/B0 , \picorv32_core/sel41_b17/B1 );
  or \picorv32_core/sel41_b17/or_B2_B3  (\picorv32_core/sel41_b17/or_B2_B3_o , \picorv32_core/sel41_b17/B2 , \picorv32_core/sel41_b17/B3 );
  or \picorv32_core/sel41_b17/or_B4_B5  (\picorv32_core/sel41_b17/or_B4_B5_o , \picorv32_core/sel41_b17/B4 , \picorv32_core/sel41_b17/B5 );
  or \picorv32_core/sel41_b17/or_B6_B7  (\picorv32_core/sel41_b17/or_B6_B7_o , \picorv32_core/sel41_b17/B6 , \picorv32_core/sel41_b17/B7 );
  or \picorv32_core/sel41_b17/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b17/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b17/or_B0_B1_o , \picorv32_core/sel41_b17/or_B2_B3_o );
  or \picorv32_core/sel41_b17/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b17/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b17/or_B4_B5_o , \picorv32_core/sel41_b17/or_B6_B7_o );
  or \picorv32_core/sel41_b17/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [17], \picorv32_core/sel41_b17/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b17/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b18/and_b0_0  (\picorv32_core/sel41_b18/B0 , \picorv32_core/n656 [18], \picorv32_core/n669 );
  and \picorv32_core/sel41_b18/and_b0_1  (\picorv32_core/sel41_b18/B1 , \picorv32_core/n584 [18], \picorv32_core/n668 );
  and \picorv32_core/sel41_b18/and_b0_2  (\picorv32_core/sel41_b18/B2 , \picorv32_core/n570 [18], \picorv32_core/n667 );
  and \picorv32_core/sel41_b18/and_b0_3  (\picorv32_core/sel41_b18/B3 , \picorv32_core/pcpi_rs1$18$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b18/and_b0_4  (\picorv32_core/sel41_b18/B4 , \picorv32_core/pcpi_rs1$18$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b18/and_b0_5  (\picorv32_core/sel41_b18/B5 , \picorv32_core/n527 [18], \picorv32_core/n664 );
  and \picorv32_core/sel41_b18/and_b0_6  (\picorv32_core/sel41_b18/B6 , \picorv32_core/pcpi_rs1$18$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b18/and_b0_7  (\picorv32_core/sel41_b18/B7 , \picorv32_core/pcpi_rs1$18$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b18/or_B0_B1  (\picorv32_core/sel41_b18/or_B0_B1_o , \picorv32_core/sel41_b18/B0 , \picorv32_core/sel41_b18/B1 );
  or \picorv32_core/sel41_b18/or_B2_B3  (\picorv32_core/sel41_b18/or_B2_B3_o , \picorv32_core/sel41_b18/B2 , \picorv32_core/sel41_b18/B3 );
  or \picorv32_core/sel41_b18/or_B4_B5  (\picorv32_core/sel41_b18/or_B4_B5_o , \picorv32_core/sel41_b18/B4 , \picorv32_core/sel41_b18/B5 );
  or \picorv32_core/sel41_b18/or_B6_B7  (\picorv32_core/sel41_b18/or_B6_B7_o , \picorv32_core/sel41_b18/B6 , \picorv32_core/sel41_b18/B7 );
  or \picorv32_core/sel41_b18/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b18/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b18/or_B0_B1_o , \picorv32_core/sel41_b18/or_B2_B3_o );
  or \picorv32_core/sel41_b18/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b18/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b18/or_B4_B5_o , \picorv32_core/sel41_b18/or_B6_B7_o );
  or \picorv32_core/sel41_b18/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [18], \picorv32_core/sel41_b18/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b18/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b19/and_b0_0  (\picorv32_core/sel41_b19/B0 , \picorv32_core/n656 [19], \picorv32_core/n669 );
  and \picorv32_core/sel41_b19/and_b0_1  (\picorv32_core/sel41_b19/B1 , \picorv32_core/n584 [19], \picorv32_core/n668 );
  and \picorv32_core/sel41_b19/and_b0_2  (\picorv32_core/sel41_b19/B2 , \picorv32_core/n570 [19], \picorv32_core/n667 );
  and \picorv32_core/sel41_b19/and_b0_3  (\picorv32_core/sel41_b19/B3 , \picorv32_core/pcpi_rs1$19$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b19/and_b0_4  (\picorv32_core/sel41_b19/B4 , \picorv32_core/pcpi_rs1$19$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b19/and_b0_5  (\picorv32_core/sel41_b19/B5 , \picorv32_core/n527 [19], \picorv32_core/n664 );
  and \picorv32_core/sel41_b19/and_b0_6  (\picorv32_core/sel41_b19/B6 , \picorv32_core/pcpi_rs1$19$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b19/and_b0_7  (\picorv32_core/sel41_b19/B7 , \picorv32_core/pcpi_rs1$19$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b19/or_B0_B1  (\picorv32_core/sel41_b19/or_B0_B1_o , \picorv32_core/sel41_b19/B0 , \picorv32_core/sel41_b19/B1 );
  or \picorv32_core/sel41_b19/or_B2_B3  (\picorv32_core/sel41_b19/or_B2_B3_o , \picorv32_core/sel41_b19/B2 , \picorv32_core/sel41_b19/B3 );
  or \picorv32_core/sel41_b19/or_B4_B5  (\picorv32_core/sel41_b19/or_B4_B5_o , \picorv32_core/sel41_b19/B4 , \picorv32_core/sel41_b19/B5 );
  or \picorv32_core/sel41_b19/or_B6_B7  (\picorv32_core/sel41_b19/or_B6_B7_o , \picorv32_core/sel41_b19/B6 , \picorv32_core/sel41_b19/B7 );
  or \picorv32_core/sel41_b19/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b19/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b19/or_B0_B1_o , \picorv32_core/sel41_b19/or_B2_B3_o );
  or \picorv32_core/sel41_b19/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b19/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b19/or_B4_B5_o , \picorv32_core/sel41_b19/or_B6_B7_o );
  or \picorv32_core/sel41_b19/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [19], \picorv32_core/sel41_b19/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b19/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b2/and_b0_0  (\picorv32_core/sel41_b2/B0 , \picorv32_core/n656 [2], \picorv32_core/n669 );
  and \picorv32_core/sel41_b2/and_b0_1  (\picorv32_core/sel41_b2/B1 , \picorv32_core/n584 [2], \picorv32_core/n668 );
  and \picorv32_core/sel41_b2/and_b0_2  (\picorv32_core/sel41_b2/B2 , \picorv32_core/n570 [2], \picorv32_core/n667 );
  and \picorv32_core/sel41_b2/and_b0_3  (\picorv32_core/sel41_b2/B3 , \picorv32_core/pcpi_rs1$2$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b2/and_b0_4  (\picorv32_core/sel41_b2/B4 , \picorv32_core/pcpi_rs1$2$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b2/and_b0_5  (\picorv32_core/sel41_b2/B5 , \picorv32_core/n527 [2], \picorv32_core/n664 );
  and \picorv32_core/sel41_b2/and_b0_6  (\picorv32_core/sel41_b2/B6 , \picorv32_core/pcpi_rs1$2$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b2/and_b0_7  (\picorv32_core/sel41_b2/B7 , \picorv32_core/pcpi_rs1$2$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b2/or_B0_B1  (\picorv32_core/sel41_b2/or_B0_B1_o , \picorv32_core/sel41_b2/B0 , \picorv32_core/sel41_b2/B1 );
  or \picorv32_core/sel41_b2/or_B2_B3  (\picorv32_core/sel41_b2/or_B2_B3_o , \picorv32_core/sel41_b2/B2 , \picorv32_core/sel41_b2/B3 );
  or \picorv32_core/sel41_b2/or_B4_B5  (\picorv32_core/sel41_b2/or_B4_B5_o , \picorv32_core/sel41_b2/B4 , \picorv32_core/sel41_b2/B5 );
  or \picorv32_core/sel41_b2/or_B6_B7  (\picorv32_core/sel41_b2/or_B6_B7_o , \picorv32_core/sel41_b2/B6 , \picorv32_core/sel41_b2/B7 );
  or \picorv32_core/sel41_b2/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b2/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b2/or_B0_B1_o , \picorv32_core/sel41_b2/or_B2_B3_o );
  or \picorv32_core/sel41_b2/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b2/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b2/or_B4_B5_o , \picorv32_core/sel41_b2/or_B6_B7_o );
  or \picorv32_core/sel41_b2/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [2], \picorv32_core/sel41_b2/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b2/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b20/and_b0_0  (\picorv32_core/sel41_b20/B0 , \picorv32_core/n656 [20], \picorv32_core/n669 );
  and \picorv32_core/sel41_b20/and_b0_1  (\picorv32_core/sel41_b20/B1 , \picorv32_core/n584 [20], \picorv32_core/n668 );
  and \picorv32_core/sel41_b20/and_b0_2  (\picorv32_core/sel41_b20/B2 , \picorv32_core/n570 [20], \picorv32_core/n667 );
  and \picorv32_core/sel41_b20/and_b0_3  (\picorv32_core/sel41_b20/B3 , \picorv32_core/pcpi_rs1$20$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b20/and_b0_4  (\picorv32_core/sel41_b20/B4 , \picorv32_core/pcpi_rs1$20$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b20/and_b0_5  (\picorv32_core/sel41_b20/B5 , \picorv32_core/n527 [20], \picorv32_core/n664 );
  and \picorv32_core/sel41_b20/and_b0_6  (\picorv32_core/sel41_b20/B6 , \picorv32_core/pcpi_rs1$20$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b20/and_b0_7  (\picorv32_core/sel41_b20/B7 , \picorv32_core/pcpi_rs1$20$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b20/or_B0_B1  (\picorv32_core/sel41_b20/or_B0_B1_o , \picorv32_core/sel41_b20/B0 , \picorv32_core/sel41_b20/B1 );
  or \picorv32_core/sel41_b20/or_B2_B3  (\picorv32_core/sel41_b20/or_B2_B3_o , \picorv32_core/sel41_b20/B2 , \picorv32_core/sel41_b20/B3 );
  or \picorv32_core/sel41_b20/or_B4_B5  (\picorv32_core/sel41_b20/or_B4_B5_o , \picorv32_core/sel41_b20/B4 , \picorv32_core/sel41_b20/B5 );
  or \picorv32_core/sel41_b20/or_B6_B7  (\picorv32_core/sel41_b20/or_B6_B7_o , \picorv32_core/sel41_b20/B6 , \picorv32_core/sel41_b20/B7 );
  or \picorv32_core/sel41_b20/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b20/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b20/or_B0_B1_o , \picorv32_core/sel41_b20/or_B2_B3_o );
  or \picorv32_core/sel41_b20/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b20/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b20/or_B4_B5_o , \picorv32_core/sel41_b20/or_B6_B7_o );
  or \picorv32_core/sel41_b20/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [20], \picorv32_core/sel41_b20/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b20/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b21/and_b0_0  (\picorv32_core/sel41_b21/B0 , \picorv32_core/n656 [21], \picorv32_core/n669 );
  and \picorv32_core/sel41_b21/and_b0_1  (\picorv32_core/sel41_b21/B1 , \picorv32_core/n584 [21], \picorv32_core/n668 );
  and \picorv32_core/sel41_b21/and_b0_2  (\picorv32_core/sel41_b21/B2 , \picorv32_core/n570 [21], \picorv32_core/n667 );
  and \picorv32_core/sel41_b21/and_b0_3  (\picorv32_core/sel41_b21/B3 , \picorv32_core/pcpi_rs1$21$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b21/and_b0_4  (\picorv32_core/sel41_b21/B4 , \picorv32_core/pcpi_rs1$21$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b21/and_b0_5  (\picorv32_core/sel41_b21/B5 , \picorv32_core/n527 [21], \picorv32_core/n664 );
  and \picorv32_core/sel41_b21/and_b0_6  (\picorv32_core/sel41_b21/B6 , \picorv32_core/pcpi_rs1$21$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b21/and_b0_7  (\picorv32_core/sel41_b21/B7 , \picorv32_core/pcpi_rs1$21$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b21/or_B0_B1  (\picorv32_core/sel41_b21/or_B0_B1_o , \picorv32_core/sel41_b21/B0 , \picorv32_core/sel41_b21/B1 );
  or \picorv32_core/sel41_b21/or_B2_B3  (\picorv32_core/sel41_b21/or_B2_B3_o , \picorv32_core/sel41_b21/B2 , \picorv32_core/sel41_b21/B3 );
  or \picorv32_core/sel41_b21/or_B4_B5  (\picorv32_core/sel41_b21/or_B4_B5_o , \picorv32_core/sel41_b21/B4 , \picorv32_core/sel41_b21/B5 );
  or \picorv32_core/sel41_b21/or_B6_B7  (\picorv32_core/sel41_b21/or_B6_B7_o , \picorv32_core/sel41_b21/B6 , \picorv32_core/sel41_b21/B7 );
  or \picorv32_core/sel41_b21/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b21/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b21/or_B0_B1_o , \picorv32_core/sel41_b21/or_B2_B3_o );
  or \picorv32_core/sel41_b21/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b21/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b21/or_B4_B5_o , \picorv32_core/sel41_b21/or_B6_B7_o );
  or \picorv32_core/sel41_b21/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [21], \picorv32_core/sel41_b21/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b21/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b22/and_b0_0  (\picorv32_core/sel41_b22/B0 , \picorv32_core/n656 [22], \picorv32_core/n669 );
  and \picorv32_core/sel41_b22/and_b0_1  (\picorv32_core/sel41_b22/B1 , \picorv32_core/n584 [22], \picorv32_core/n668 );
  and \picorv32_core/sel41_b22/and_b0_2  (\picorv32_core/sel41_b22/B2 , \picorv32_core/n570 [22], \picorv32_core/n667 );
  and \picorv32_core/sel41_b22/and_b0_3  (\picorv32_core/sel41_b22/B3 , \picorv32_core/pcpi_rs1$22$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b22/and_b0_4  (\picorv32_core/sel41_b22/B4 , \picorv32_core/pcpi_rs1$22$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b22/and_b0_5  (\picorv32_core/sel41_b22/B5 , \picorv32_core/n527 [22], \picorv32_core/n664 );
  and \picorv32_core/sel41_b22/and_b0_6  (\picorv32_core/sel41_b22/B6 , \picorv32_core/pcpi_rs1$22$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b22/and_b0_7  (\picorv32_core/sel41_b22/B7 , \picorv32_core/pcpi_rs1$22$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b22/or_B0_B1  (\picorv32_core/sel41_b22/or_B0_B1_o , \picorv32_core/sel41_b22/B0 , \picorv32_core/sel41_b22/B1 );
  or \picorv32_core/sel41_b22/or_B2_B3  (\picorv32_core/sel41_b22/or_B2_B3_o , \picorv32_core/sel41_b22/B2 , \picorv32_core/sel41_b22/B3 );
  or \picorv32_core/sel41_b22/or_B4_B5  (\picorv32_core/sel41_b22/or_B4_B5_o , \picorv32_core/sel41_b22/B4 , \picorv32_core/sel41_b22/B5 );
  or \picorv32_core/sel41_b22/or_B6_B7  (\picorv32_core/sel41_b22/or_B6_B7_o , \picorv32_core/sel41_b22/B6 , \picorv32_core/sel41_b22/B7 );
  or \picorv32_core/sel41_b22/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b22/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b22/or_B0_B1_o , \picorv32_core/sel41_b22/or_B2_B3_o );
  or \picorv32_core/sel41_b22/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b22/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b22/or_B4_B5_o , \picorv32_core/sel41_b22/or_B6_B7_o );
  or \picorv32_core/sel41_b22/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [22], \picorv32_core/sel41_b22/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b22/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b23/and_b0_0  (\picorv32_core/sel41_b23/B0 , \picorv32_core/n656 [23], \picorv32_core/n669 );
  and \picorv32_core/sel41_b23/and_b0_1  (\picorv32_core/sel41_b23/B1 , \picorv32_core/n584 [23], \picorv32_core/n668 );
  and \picorv32_core/sel41_b23/and_b0_2  (\picorv32_core/sel41_b23/B2 , \picorv32_core/n570 [23], \picorv32_core/n667 );
  and \picorv32_core/sel41_b23/and_b0_3  (\picorv32_core/sel41_b23/B3 , \picorv32_core/pcpi_rs1$23$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b23/and_b0_4  (\picorv32_core/sel41_b23/B4 , \picorv32_core/pcpi_rs1$23$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b23/and_b0_5  (\picorv32_core/sel41_b23/B5 , \picorv32_core/n527 [23], \picorv32_core/n664 );
  and \picorv32_core/sel41_b23/and_b0_6  (\picorv32_core/sel41_b23/B6 , \picorv32_core/pcpi_rs1$23$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b23/and_b0_7  (\picorv32_core/sel41_b23/B7 , \picorv32_core/pcpi_rs1$23$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b23/or_B0_B1  (\picorv32_core/sel41_b23/or_B0_B1_o , \picorv32_core/sel41_b23/B0 , \picorv32_core/sel41_b23/B1 );
  or \picorv32_core/sel41_b23/or_B2_B3  (\picorv32_core/sel41_b23/or_B2_B3_o , \picorv32_core/sel41_b23/B2 , \picorv32_core/sel41_b23/B3 );
  or \picorv32_core/sel41_b23/or_B4_B5  (\picorv32_core/sel41_b23/or_B4_B5_o , \picorv32_core/sel41_b23/B4 , \picorv32_core/sel41_b23/B5 );
  or \picorv32_core/sel41_b23/or_B6_B7  (\picorv32_core/sel41_b23/or_B6_B7_o , \picorv32_core/sel41_b23/B6 , \picorv32_core/sel41_b23/B7 );
  or \picorv32_core/sel41_b23/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b23/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b23/or_B0_B1_o , \picorv32_core/sel41_b23/or_B2_B3_o );
  or \picorv32_core/sel41_b23/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b23/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b23/or_B4_B5_o , \picorv32_core/sel41_b23/or_B6_B7_o );
  or \picorv32_core/sel41_b23/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [23], \picorv32_core/sel41_b23/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b23/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b24/and_b0_0  (\picorv32_core/sel41_b24/B0 , \picorv32_core/n656 [24], \picorv32_core/n669 );
  and \picorv32_core/sel41_b24/and_b0_1  (\picorv32_core/sel41_b24/B1 , \picorv32_core/n584 [24], \picorv32_core/n668 );
  and \picorv32_core/sel41_b24/and_b0_2  (\picorv32_core/sel41_b24/B2 , \picorv32_core/n570 [24], \picorv32_core/n667 );
  and \picorv32_core/sel41_b24/and_b0_3  (\picorv32_core/sel41_b24/B3 , \picorv32_core/pcpi_rs1$24$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b24/and_b0_4  (\picorv32_core/sel41_b24/B4 , \picorv32_core/pcpi_rs1$24$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b24/and_b0_5  (\picorv32_core/sel41_b24/B5 , \picorv32_core/n527 [24], \picorv32_core/n664 );
  and \picorv32_core/sel41_b24/and_b0_6  (\picorv32_core/sel41_b24/B6 , \picorv32_core/pcpi_rs1$24$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b24/and_b0_7  (\picorv32_core/sel41_b24/B7 , \picorv32_core/pcpi_rs1$24$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b24/or_B0_B1  (\picorv32_core/sel41_b24/or_B0_B1_o , \picorv32_core/sel41_b24/B0 , \picorv32_core/sel41_b24/B1 );
  or \picorv32_core/sel41_b24/or_B2_B3  (\picorv32_core/sel41_b24/or_B2_B3_o , \picorv32_core/sel41_b24/B2 , \picorv32_core/sel41_b24/B3 );
  or \picorv32_core/sel41_b24/or_B4_B5  (\picorv32_core/sel41_b24/or_B4_B5_o , \picorv32_core/sel41_b24/B4 , \picorv32_core/sel41_b24/B5 );
  or \picorv32_core/sel41_b24/or_B6_B7  (\picorv32_core/sel41_b24/or_B6_B7_o , \picorv32_core/sel41_b24/B6 , \picorv32_core/sel41_b24/B7 );
  or \picorv32_core/sel41_b24/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b24/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b24/or_B0_B1_o , \picorv32_core/sel41_b24/or_B2_B3_o );
  or \picorv32_core/sel41_b24/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b24/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b24/or_B4_B5_o , \picorv32_core/sel41_b24/or_B6_B7_o );
  or \picorv32_core/sel41_b24/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [24], \picorv32_core/sel41_b24/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b24/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b25/and_b0_0  (\picorv32_core/sel41_b25/B0 , \picorv32_core/n656 [25], \picorv32_core/n669 );
  and \picorv32_core/sel41_b25/and_b0_1  (\picorv32_core/sel41_b25/B1 , \picorv32_core/n584 [25], \picorv32_core/n668 );
  and \picorv32_core/sel41_b25/and_b0_2  (\picorv32_core/sel41_b25/B2 , \picorv32_core/n570 [25], \picorv32_core/n667 );
  and \picorv32_core/sel41_b25/and_b0_3  (\picorv32_core/sel41_b25/B3 , \picorv32_core/pcpi_rs1$25$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b25/and_b0_4  (\picorv32_core/sel41_b25/B4 , \picorv32_core/pcpi_rs1$25$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b25/and_b0_5  (\picorv32_core/sel41_b25/B5 , \picorv32_core/n527 [25], \picorv32_core/n664 );
  and \picorv32_core/sel41_b25/and_b0_6  (\picorv32_core/sel41_b25/B6 , \picorv32_core/pcpi_rs1$25$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b25/and_b0_7  (\picorv32_core/sel41_b25/B7 , \picorv32_core/pcpi_rs1$25$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b25/or_B0_B1  (\picorv32_core/sel41_b25/or_B0_B1_o , \picorv32_core/sel41_b25/B0 , \picorv32_core/sel41_b25/B1 );
  or \picorv32_core/sel41_b25/or_B2_B3  (\picorv32_core/sel41_b25/or_B2_B3_o , \picorv32_core/sel41_b25/B2 , \picorv32_core/sel41_b25/B3 );
  or \picorv32_core/sel41_b25/or_B4_B5  (\picorv32_core/sel41_b25/or_B4_B5_o , \picorv32_core/sel41_b25/B4 , \picorv32_core/sel41_b25/B5 );
  or \picorv32_core/sel41_b25/or_B6_B7  (\picorv32_core/sel41_b25/or_B6_B7_o , \picorv32_core/sel41_b25/B6 , \picorv32_core/sel41_b25/B7 );
  or \picorv32_core/sel41_b25/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b25/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b25/or_B0_B1_o , \picorv32_core/sel41_b25/or_B2_B3_o );
  or \picorv32_core/sel41_b25/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b25/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b25/or_B4_B5_o , \picorv32_core/sel41_b25/or_B6_B7_o );
  or \picorv32_core/sel41_b25/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [25], \picorv32_core/sel41_b25/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b25/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b26/and_b0_0  (\picorv32_core/sel41_b26/B0 , \picorv32_core/n656 [26], \picorv32_core/n669 );
  and \picorv32_core/sel41_b26/and_b0_1  (\picorv32_core/sel41_b26/B1 , \picorv32_core/n584 [26], \picorv32_core/n668 );
  and \picorv32_core/sel41_b26/and_b0_2  (\picorv32_core/sel41_b26/B2 , \picorv32_core/n570 [26], \picorv32_core/n667 );
  and \picorv32_core/sel41_b26/and_b0_3  (\picorv32_core/sel41_b26/B3 , \picorv32_core/pcpi_rs1$26$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b26/and_b0_4  (\picorv32_core/sel41_b26/B4 , \picorv32_core/pcpi_rs1$26$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b26/and_b0_5  (\picorv32_core/sel41_b26/B5 , \picorv32_core/n527 [26], \picorv32_core/n664 );
  and \picorv32_core/sel41_b26/and_b0_6  (\picorv32_core/sel41_b26/B6 , \picorv32_core/pcpi_rs1$26$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b26/and_b0_7  (\picorv32_core/sel41_b26/B7 , \picorv32_core/pcpi_rs1$26$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b26/or_B0_B1  (\picorv32_core/sel41_b26/or_B0_B1_o , \picorv32_core/sel41_b26/B0 , \picorv32_core/sel41_b26/B1 );
  or \picorv32_core/sel41_b26/or_B2_B3  (\picorv32_core/sel41_b26/or_B2_B3_o , \picorv32_core/sel41_b26/B2 , \picorv32_core/sel41_b26/B3 );
  or \picorv32_core/sel41_b26/or_B4_B5  (\picorv32_core/sel41_b26/or_B4_B5_o , \picorv32_core/sel41_b26/B4 , \picorv32_core/sel41_b26/B5 );
  or \picorv32_core/sel41_b26/or_B6_B7  (\picorv32_core/sel41_b26/or_B6_B7_o , \picorv32_core/sel41_b26/B6 , \picorv32_core/sel41_b26/B7 );
  or \picorv32_core/sel41_b26/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b26/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b26/or_B0_B1_o , \picorv32_core/sel41_b26/or_B2_B3_o );
  or \picorv32_core/sel41_b26/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b26/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b26/or_B4_B5_o , \picorv32_core/sel41_b26/or_B6_B7_o );
  or \picorv32_core/sel41_b26/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [26], \picorv32_core/sel41_b26/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b26/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b27/and_b0_0  (\picorv32_core/sel41_b27/B0 , \picorv32_core/n656 [27], \picorv32_core/n669 );
  and \picorv32_core/sel41_b27/and_b0_1  (\picorv32_core/sel41_b27/B1 , \picorv32_core/n584 [27], \picorv32_core/n668 );
  and \picorv32_core/sel41_b27/and_b0_2  (\picorv32_core/sel41_b27/B2 , \picorv32_core/n570 [27], \picorv32_core/n667 );
  and \picorv32_core/sel41_b27/and_b0_3  (\picorv32_core/sel41_b27/B3 , \picorv32_core/pcpi_rs1$27$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b27/and_b0_4  (\picorv32_core/sel41_b27/B4 , \picorv32_core/pcpi_rs1$27$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b27/and_b0_5  (\picorv32_core/sel41_b27/B5 , \picorv32_core/n527 [27], \picorv32_core/n664 );
  and \picorv32_core/sel41_b27/and_b0_6  (\picorv32_core/sel41_b27/B6 , \picorv32_core/pcpi_rs1$27$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b27/and_b0_7  (\picorv32_core/sel41_b27/B7 , \picorv32_core/pcpi_rs1$27$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b27/or_B0_B1  (\picorv32_core/sel41_b27/or_B0_B1_o , \picorv32_core/sel41_b27/B0 , \picorv32_core/sel41_b27/B1 );
  or \picorv32_core/sel41_b27/or_B2_B3  (\picorv32_core/sel41_b27/or_B2_B3_o , \picorv32_core/sel41_b27/B2 , \picorv32_core/sel41_b27/B3 );
  or \picorv32_core/sel41_b27/or_B4_B5  (\picorv32_core/sel41_b27/or_B4_B5_o , \picorv32_core/sel41_b27/B4 , \picorv32_core/sel41_b27/B5 );
  or \picorv32_core/sel41_b27/or_B6_B7  (\picorv32_core/sel41_b27/or_B6_B7_o , \picorv32_core/sel41_b27/B6 , \picorv32_core/sel41_b27/B7 );
  or \picorv32_core/sel41_b27/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b27/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b27/or_B0_B1_o , \picorv32_core/sel41_b27/or_B2_B3_o );
  or \picorv32_core/sel41_b27/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b27/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b27/or_B4_B5_o , \picorv32_core/sel41_b27/or_B6_B7_o );
  or \picorv32_core/sel41_b27/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [27], \picorv32_core/sel41_b27/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b27/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b28/and_b0_0  (\picorv32_core/sel41_b28/B0 , \picorv32_core/n656 [28], \picorv32_core/n669 );
  and \picorv32_core/sel41_b28/and_b0_1  (\picorv32_core/sel41_b28/B1 , \picorv32_core/n584 [28], \picorv32_core/n668 );
  and \picorv32_core/sel41_b28/and_b0_2  (\picorv32_core/sel41_b28/B2 , \picorv32_core/n570 [28], \picorv32_core/n667 );
  and \picorv32_core/sel41_b28/and_b0_3  (\picorv32_core/sel41_b28/B3 , \picorv32_core/pcpi_rs1$28$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b28/and_b0_4  (\picorv32_core/sel41_b28/B4 , \picorv32_core/pcpi_rs1$28$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b28/and_b0_5  (\picorv32_core/sel41_b28/B5 , \picorv32_core/n527 [28], \picorv32_core/n664 );
  and \picorv32_core/sel41_b28/and_b0_6  (\picorv32_core/sel41_b28/B6 , \picorv32_core/pcpi_rs1$28$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b28/and_b0_7  (\picorv32_core/sel41_b28/B7 , \picorv32_core/pcpi_rs1$28$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b28/or_B0_B1  (\picorv32_core/sel41_b28/or_B0_B1_o , \picorv32_core/sel41_b28/B0 , \picorv32_core/sel41_b28/B1 );
  or \picorv32_core/sel41_b28/or_B2_B3  (\picorv32_core/sel41_b28/or_B2_B3_o , \picorv32_core/sel41_b28/B2 , \picorv32_core/sel41_b28/B3 );
  or \picorv32_core/sel41_b28/or_B4_B5  (\picorv32_core/sel41_b28/or_B4_B5_o , \picorv32_core/sel41_b28/B4 , \picorv32_core/sel41_b28/B5 );
  or \picorv32_core/sel41_b28/or_B6_B7  (\picorv32_core/sel41_b28/or_B6_B7_o , \picorv32_core/sel41_b28/B6 , \picorv32_core/sel41_b28/B7 );
  or \picorv32_core/sel41_b28/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b28/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b28/or_B0_B1_o , \picorv32_core/sel41_b28/or_B2_B3_o );
  or \picorv32_core/sel41_b28/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b28/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b28/or_B4_B5_o , \picorv32_core/sel41_b28/or_B6_B7_o );
  or \picorv32_core/sel41_b28/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [28], \picorv32_core/sel41_b28/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b28/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b29/and_b0_0  (\picorv32_core/sel41_b29/B0 , \picorv32_core/n656 [29], \picorv32_core/n669 );
  and \picorv32_core/sel41_b29/and_b0_1  (\picorv32_core/sel41_b29/B1 , \picorv32_core/n584 [29], \picorv32_core/n668 );
  and \picorv32_core/sel41_b29/and_b0_2  (\picorv32_core/sel41_b29/B2 , \picorv32_core/n570 [29], \picorv32_core/n667 );
  and \picorv32_core/sel41_b29/and_b0_3  (\picorv32_core/sel41_b29/B3 , \picorv32_core/pcpi_rs1$29$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b29/and_b0_4  (\picorv32_core/sel41_b29/B4 , \picorv32_core/pcpi_rs1$29$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b29/and_b0_5  (\picorv32_core/sel41_b29/B5 , \picorv32_core/n527 [29], \picorv32_core/n664 );
  and \picorv32_core/sel41_b29/and_b0_6  (\picorv32_core/sel41_b29/B6 , \picorv32_core/pcpi_rs1$29$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b29/and_b0_7  (\picorv32_core/sel41_b29/B7 , \picorv32_core/pcpi_rs1$29$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b29/or_B0_B1  (\picorv32_core/sel41_b29/or_B0_B1_o , \picorv32_core/sel41_b29/B0 , \picorv32_core/sel41_b29/B1 );
  or \picorv32_core/sel41_b29/or_B2_B3  (\picorv32_core/sel41_b29/or_B2_B3_o , \picorv32_core/sel41_b29/B2 , \picorv32_core/sel41_b29/B3 );
  or \picorv32_core/sel41_b29/or_B4_B5  (\picorv32_core/sel41_b29/or_B4_B5_o , \picorv32_core/sel41_b29/B4 , \picorv32_core/sel41_b29/B5 );
  or \picorv32_core/sel41_b29/or_B6_B7  (\picorv32_core/sel41_b29/or_B6_B7_o , \picorv32_core/sel41_b29/B6 , \picorv32_core/sel41_b29/B7 );
  or \picorv32_core/sel41_b29/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b29/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b29/or_B0_B1_o , \picorv32_core/sel41_b29/or_B2_B3_o );
  or \picorv32_core/sel41_b29/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b29/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b29/or_B4_B5_o , \picorv32_core/sel41_b29/or_B6_B7_o );
  or \picorv32_core/sel41_b29/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [29], \picorv32_core/sel41_b29/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b29/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b3/and_b0_0  (\picorv32_core/sel41_b3/B0 , \picorv32_core/n656 [3], \picorv32_core/n669 );
  and \picorv32_core/sel41_b3/and_b0_1  (\picorv32_core/sel41_b3/B1 , \picorv32_core/n584 [3], \picorv32_core/n668 );
  and \picorv32_core/sel41_b3/and_b0_2  (\picorv32_core/sel41_b3/B2 , \picorv32_core/n570 [3], \picorv32_core/n667 );
  and \picorv32_core/sel41_b3/and_b0_3  (\picorv32_core/sel41_b3/B3 , \picorv32_core/pcpi_rs1$3$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b3/and_b0_4  (\picorv32_core/sel41_b3/B4 , \picorv32_core/pcpi_rs1$3$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b3/and_b0_5  (\picorv32_core/sel41_b3/B5 , \picorv32_core/n527 [3], \picorv32_core/n664 );
  and \picorv32_core/sel41_b3/and_b0_6  (\picorv32_core/sel41_b3/B6 , \picorv32_core/pcpi_rs1$3$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b3/and_b0_7  (\picorv32_core/sel41_b3/B7 , \picorv32_core/pcpi_rs1$3$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b3/or_B0_B1  (\picorv32_core/sel41_b3/or_B0_B1_o , \picorv32_core/sel41_b3/B0 , \picorv32_core/sel41_b3/B1 );
  or \picorv32_core/sel41_b3/or_B2_B3  (\picorv32_core/sel41_b3/or_B2_B3_o , \picorv32_core/sel41_b3/B2 , \picorv32_core/sel41_b3/B3 );
  or \picorv32_core/sel41_b3/or_B4_B5  (\picorv32_core/sel41_b3/or_B4_B5_o , \picorv32_core/sel41_b3/B4 , \picorv32_core/sel41_b3/B5 );
  or \picorv32_core/sel41_b3/or_B6_B7  (\picorv32_core/sel41_b3/or_B6_B7_o , \picorv32_core/sel41_b3/B6 , \picorv32_core/sel41_b3/B7 );
  or \picorv32_core/sel41_b3/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b3/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b3/or_B0_B1_o , \picorv32_core/sel41_b3/or_B2_B3_o );
  or \picorv32_core/sel41_b3/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b3/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b3/or_B4_B5_o , \picorv32_core/sel41_b3/or_B6_B7_o );
  or \picorv32_core/sel41_b3/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [3], \picorv32_core/sel41_b3/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b3/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b30/and_b0_0  (\picorv32_core/sel41_b30/B0 , \picorv32_core/n656 [30], \picorv32_core/n669 );
  and \picorv32_core/sel41_b30/and_b0_1  (\picorv32_core/sel41_b30/B1 , \picorv32_core/n584 [30], \picorv32_core/n668 );
  and \picorv32_core/sel41_b30/and_b0_2  (\picorv32_core/sel41_b30/B2 , \picorv32_core/n570 [30], \picorv32_core/n667 );
  and \picorv32_core/sel41_b30/and_b0_3  (\picorv32_core/sel41_b30/B3 , \picorv32_core/pcpi_rs1$30$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b30/and_b0_4  (\picorv32_core/sel41_b30/B4 , \picorv32_core/pcpi_rs1$30$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b30/and_b0_5  (\picorv32_core/sel41_b30/B5 , \picorv32_core/n527 [30], \picorv32_core/n664 );
  and \picorv32_core/sel41_b30/and_b0_6  (\picorv32_core/sel41_b30/B6 , \picorv32_core/pcpi_rs1$30$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b30/and_b0_7  (\picorv32_core/sel41_b30/B7 , \picorv32_core/pcpi_rs1$30$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b30/or_B0_B1  (\picorv32_core/sel41_b30/or_B0_B1_o , \picorv32_core/sel41_b30/B0 , \picorv32_core/sel41_b30/B1 );
  or \picorv32_core/sel41_b30/or_B2_B3  (\picorv32_core/sel41_b30/or_B2_B3_o , \picorv32_core/sel41_b30/B2 , \picorv32_core/sel41_b30/B3 );
  or \picorv32_core/sel41_b30/or_B4_B5  (\picorv32_core/sel41_b30/or_B4_B5_o , \picorv32_core/sel41_b30/B4 , \picorv32_core/sel41_b30/B5 );
  or \picorv32_core/sel41_b30/or_B6_B7  (\picorv32_core/sel41_b30/or_B6_B7_o , \picorv32_core/sel41_b30/B6 , \picorv32_core/sel41_b30/B7 );
  or \picorv32_core/sel41_b30/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b30/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b30/or_B0_B1_o , \picorv32_core/sel41_b30/or_B2_B3_o );
  or \picorv32_core/sel41_b30/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b30/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b30/or_B4_B5_o , \picorv32_core/sel41_b30/or_B6_B7_o );
  or \picorv32_core/sel41_b30/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [30], \picorv32_core/sel41_b30/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b30/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b31/and_b0_0  (\picorv32_core/sel41_b31/B0 , \picorv32_core/n656 [31], \picorv32_core/n669 );
  and \picorv32_core/sel41_b31/and_b0_1  (\picorv32_core/sel41_b31/B1 , \picorv32_core/n584 [31], \picorv32_core/n668 );
  and \picorv32_core/sel41_b31/and_b0_2  (\picorv32_core/sel41_b31/B2 , \picorv32_core/n570 [31], \picorv32_core/n667 );
  and \picorv32_core/sel41_b31/and_b0_3  (\picorv32_core/sel41_b31/B3 , \picorv32_core/pcpi_rs1$31$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b31/and_b0_4  (\picorv32_core/sel41_b31/B4 , \picorv32_core/pcpi_rs1$31$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b31/and_b0_5  (\picorv32_core/sel41_b31/B5 , \picorv32_core/n527 [31], \picorv32_core/n664 );
  and \picorv32_core/sel41_b31/and_b0_6  (\picorv32_core/sel41_b31/B6 , \picorv32_core/pcpi_rs1$31$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b31/and_b0_7  (\picorv32_core/sel41_b31/B7 , \picorv32_core/pcpi_rs1$31$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b31/or_B0_B1  (\picorv32_core/sel41_b31/or_B0_B1_o , \picorv32_core/sel41_b31/B0 , \picorv32_core/sel41_b31/B1 );
  or \picorv32_core/sel41_b31/or_B2_B3  (\picorv32_core/sel41_b31/or_B2_B3_o , \picorv32_core/sel41_b31/B2 , \picorv32_core/sel41_b31/B3 );
  or \picorv32_core/sel41_b31/or_B4_B5  (\picorv32_core/sel41_b31/or_B4_B5_o , \picorv32_core/sel41_b31/B4 , \picorv32_core/sel41_b31/B5 );
  or \picorv32_core/sel41_b31/or_B6_B7  (\picorv32_core/sel41_b31/or_B6_B7_o , \picorv32_core/sel41_b31/B6 , \picorv32_core/sel41_b31/B7 );
  or \picorv32_core/sel41_b31/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b31/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b31/or_B0_B1_o , \picorv32_core/sel41_b31/or_B2_B3_o );
  or \picorv32_core/sel41_b31/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b31/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b31/or_B4_B5_o , \picorv32_core/sel41_b31/or_B6_B7_o );
  or \picorv32_core/sel41_b31/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [31], \picorv32_core/sel41_b31/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b31/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b4/and_b0_0  (\picorv32_core/sel41_b4/B0 , \picorv32_core/n656 [4], \picorv32_core/n669 );
  and \picorv32_core/sel41_b4/and_b0_1  (\picorv32_core/sel41_b4/B1 , \picorv32_core/n584 [4], \picorv32_core/n668 );
  and \picorv32_core/sel41_b4/and_b0_2  (\picorv32_core/sel41_b4/B2 , \picorv32_core/n570 [4], \picorv32_core/n667 );
  and \picorv32_core/sel41_b4/and_b0_3  (\picorv32_core/sel41_b4/B3 , \picorv32_core/pcpi_rs1$4$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b4/and_b0_4  (\picorv32_core/sel41_b4/B4 , \picorv32_core/pcpi_rs1$4$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b4/and_b0_5  (\picorv32_core/sel41_b4/B5 , \picorv32_core/n527 [4], \picorv32_core/n664 );
  and \picorv32_core/sel41_b4/and_b0_6  (\picorv32_core/sel41_b4/B6 , \picorv32_core/pcpi_rs1$4$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b4/and_b0_7  (\picorv32_core/sel41_b4/B7 , \picorv32_core/pcpi_rs1$4$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b4/or_B0_B1  (\picorv32_core/sel41_b4/or_B0_B1_o , \picorv32_core/sel41_b4/B0 , \picorv32_core/sel41_b4/B1 );
  or \picorv32_core/sel41_b4/or_B2_B3  (\picorv32_core/sel41_b4/or_B2_B3_o , \picorv32_core/sel41_b4/B2 , \picorv32_core/sel41_b4/B3 );
  or \picorv32_core/sel41_b4/or_B4_B5  (\picorv32_core/sel41_b4/or_B4_B5_o , \picorv32_core/sel41_b4/B4 , \picorv32_core/sel41_b4/B5 );
  or \picorv32_core/sel41_b4/or_B6_B7  (\picorv32_core/sel41_b4/or_B6_B7_o , \picorv32_core/sel41_b4/B6 , \picorv32_core/sel41_b4/B7 );
  or \picorv32_core/sel41_b4/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b4/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b4/or_B0_B1_o , \picorv32_core/sel41_b4/or_B2_B3_o );
  or \picorv32_core/sel41_b4/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b4/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b4/or_B4_B5_o , \picorv32_core/sel41_b4/or_B6_B7_o );
  or \picorv32_core/sel41_b4/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [4], \picorv32_core/sel41_b4/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b4/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b5/and_b0_0  (\picorv32_core/sel41_b5/B0 , \picorv32_core/n656 [5], \picorv32_core/n669 );
  and \picorv32_core/sel41_b5/and_b0_1  (\picorv32_core/sel41_b5/B1 , \picorv32_core/n584 [5], \picorv32_core/n668 );
  and \picorv32_core/sel41_b5/and_b0_2  (\picorv32_core/sel41_b5/B2 , \picorv32_core/n570 [5], \picorv32_core/n667 );
  and \picorv32_core/sel41_b5/and_b0_3  (\picorv32_core/sel41_b5/B3 , \picorv32_core/pcpi_rs1$5$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b5/and_b0_4  (\picorv32_core/sel41_b5/B4 , \picorv32_core/pcpi_rs1$5$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b5/and_b0_5  (\picorv32_core/sel41_b5/B5 , \picorv32_core/n527 [5], \picorv32_core/n664 );
  and \picorv32_core/sel41_b5/and_b0_6  (\picorv32_core/sel41_b5/B6 , \picorv32_core/pcpi_rs1$5$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b5/and_b0_7  (\picorv32_core/sel41_b5/B7 , \picorv32_core/pcpi_rs1$5$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b5/or_B0_B1  (\picorv32_core/sel41_b5/or_B0_B1_o , \picorv32_core/sel41_b5/B0 , \picorv32_core/sel41_b5/B1 );
  or \picorv32_core/sel41_b5/or_B2_B3  (\picorv32_core/sel41_b5/or_B2_B3_o , \picorv32_core/sel41_b5/B2 , \picorv32_core/sel41_b5/B3 );
  or \picorv32_core/sel41_b5/or_B4_B5  (\picorv32_core/sel41_b5/or_B4_B5_o , \picorv32_core/sel41_b5/B4 , \picorv32_core/sel41_b5/B5 );
  or \picorv32_core/sel41_b5/or_B6_B7  (\picorv32_core/sel41_b5/or_B6_B7_o , \picorv32_core/sel41_b5/B6 , \picorv32_core/sel41_b5/B7 );
  or \picorv32_core/sel41_b5/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b5/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b5/or_B0_B1_o , \picorv32_core/sel41_b5/or_B2_B3_o );
  or \picorv32_core/sel41_b5/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b5/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b5/or_B4_B5_o , \picorv32_core/sel41_b5/or_B6_B7_o );
  or \picorv32_core/sel41_b5/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [5], \picorv32_core/sel41_b5/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b5/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b6/and_b0_0  (\picorv32_core/sel41_b6/B0 , \picorv32_core/n656 [6], \picorv32_core/n669 );
  and \picorv32_core/sel41_b6/and_b0_1  (\picorv32_core/sel41_b6/B1 , \picorv32_core/n584 [6], \picorv32_core/n668 );
  and \picorv32_core/sel41_b6/and_b0_2  (\picorv32_core/sel41_b6/B2 , \picorv32_core/n570 [6], \picorv32_core/n667 );
  and \picorv32_core/sel41_b6/and_b0_3  (\picorv32_core/sel41_b6/B3 , \picorv32_core/pcpi_rs1$6$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b6/and_b0_4  (\picorv32_core/sel41_b6/B4 , \picorv32_core/pcpi_rs1$6$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b6/and_b0_5  (\picorv32_core/sel41_b6/B5 , \picorv32_core/n527 [6], \picorv32_core/n664 );
  and \picorv32_core/sel41_b6/and_b0_6  (\picorv32_core/sel41_b6/B6 , \picorv32_core/pcpi_rs1$6$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b6/and_b0_7  (\picorv32_core/sel41_b6/B7 , \picorv32_core/pcpi_rs1$6$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b6/or_B0_B1  (\picorv32_core/sel41_b6/or_B0_B1_o , \picorv32_core/sel41_b6/B0 , \picorv32_core/sel41_b6/B1 );
  or \picorv32_core/sel41_b6/or_B2_B3  (\picorv32_core/sel41_b6/or_B2_B3_o , \picorv32_core/sel41_b6/B2 , \picorv32_core/sel41_b6/B3 );
  or \picorv32_core/sel41_b6/or_B4_B5  (\picorv32_core/sel41_b6/or_B4_B5_o , \picorv32_core/sel41_b6/B4 , \picorv32_core/sel41_b6/B5 );
  or \picorv32_core/sel41_b6/or_B6_B7  (\picorv32_core/sel41_b6/or_B6_B7_o , \picorv32_core/sel41_b6/B6 , \picorv32_core/sel41_b6/B7 );
  or \picorv32_core/sel41_b6/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b6/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b6/or_B0_B1_o , \picorv32_core/sel41_b6/or_B2_B3_o );
  or \picorv32_core/sel41_b6/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b6/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b6/or_B4_B5_o , \picorv32_core/sel41_b6/or_B6_B7_o );
  or \picorv32_core/sel41_b6/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [6], \picorv32_core/sel41_b6/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b6/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b7/and_b0_0  (\picorv32_core/sel41_b7/B0 , \picorv32_core/n656 [7], \picorv32_core/n669 );
  and \picorv32_core/sel41_b7/and_b0_1  (\picorv32_core/sel41_b7/B1 , \picorv32_core/n584 [7], \picorv32_core/n668 );
  and \picorv32_core/sel41_b7/and_b0_2  (\picorv32_core/sel41_b7/B2 , \picorv32_core/n570 [7], \picorv32_core/n667 );
  and \picorv32_core/sel41_b7/and_b0_3  (\picorv32_core/sel41_b7/B3 , \picorv32_core/pcpi_rs1$7$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b7/and_b0_4  (\picorv32_core/sel41_b7/B4 , \picorv32_core/pcpi_rs1$7$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b7/and_b0_5  (\picorv32_core/sel41_b7/B5 , \picorv32_core/n527 [7], \picorv32_core/n664 );
  and \picorv32_core/sel41_b7/and_b0_6  (\picorv32_core/sel41_b7/B6 , \picorv32_core/pcpi_rs1$7$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b7/and_b0_7  (\picorv32_core/sel41_b7/B7 , \picorv32_core/pcpi_rs1$7$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b7/or_B0_B1  (\picorv32_core/sel41_b7/or_B0_B1_o , \picorv32_core/sel41_b7/B0 , \picorv32_core/sel41_b7/B1 );
  or \picorv32_core/sel41_b7/or_B2_B3  (\picorv32_core/sel41_b7/or_B2_B3_o , \picorv32_core/sel41_b7/B2 , \picorv32_core/sel41_b7/B3 );
  or \picorv32_core/sel41_b7/or_B4_B5  (\picorv32_core/sel41_b7/or_B4_B5_o , \picorv32_core/sel41_b7/B4 , \picorv32_core/sel41_b7/B5 );
  or \picorv32_core/sel41_b7/or_B6_B7  (\picorv32_core/sel41_b7/or_B6_B7_o , \picorv32_core/sel41_b7/B6 , \picorv32_core/sel41_b7/B7 );
  or \picorv32_core/sel41_b7/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b7/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b7/or_B0_B1_o , \picorv32_core/sel41_b7/or_B2_B3_o );
  or \picorv32_core/sel41_b7/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b7/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b7/or_B4_B5_o , \picorv32_core/sel41_b7/or_B6_B7_o );
  or \picorv32_core/sel41_b7/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [7], \picorv32_core/sel41_b7/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b7/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b8/and_b0_0  (\picorv32_core/sel41_b8/B0 , \picorv32_core/n656 [8], \picorv32_core/n669 );
  and \picorv32_core/sel41_b8/and_b0_1  (\picorv32_core/sel41_b8/B1 , \picorv32_core/n584 [8], \picorv32_core/n668 );
  and \picorv32_core/sel41_b8/and_b0_2  (\picorv32_core/sel41_b8/B2 , \picorv32_core/n570 [8], \picorv32_core/n667 );
  and \picorv32_core/sel41_b8/and_b0_3  (\picorv32_core/sel41_b8/B3 , \picorv32_core/pcpi_rs1$8$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b8/and_b0_4  (\picorv32_core/sel41_b8/B4 , \picorv32_core/pcpi_rs1$8$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b8/and_b0_5  (\picorv32_core/sel41_b8/B5 , \picorv32_core/n527 [8], \picorv32_core/n664 );
  and \picorv32_core/sel41_b8/and_b0_6  (\picorv32_core/sel41_b8/B6 , \picorv32_core/pcpi_rs1$8$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b8/and_b0_7  (\picorv32_core/sel41_b8/B7 , \picorv32_core/pcpi_rs1$8$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b8/or_B0_B1  (\picorv32_core/sel41_b8/or_B0_B1_o , \picorv32_core/sel41_b8/B0 , \picorv32_core/sel41_b8/B1 );
  or \picorv32_core/sel41_b8/or_B2_B3  (\picorv32_core/sel41_b8/or_B2_B3_o , \picorv32_core/sel41_b8/B2 , \picorv32_core/sel41_b8/B3 );
  or \picorv32_core/sel41_b8/or_B4_B5  (\picorv32_core/sel41_b8/or_B4_B5_o , \picorv32_core/sel41_b8/B4 , \picorv32_core/sel41_b8/B5 );
  or \picorv32_core/sel41_b8/or_B6_B7  (\picorv32_core/sel41_b8/or_B6_B7_o , \picorv32_core/sel41_b8/B6 , \picorv32_core/sel41_b8/B7 );
  or \picorv32_core/sel41_b8/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b8/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b8/or_B0_B1_o , \picorv32_core/sel41_b8/or_B2_B3_o );
  or \picorv32_core/sel41_b8/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b8/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b8/or_B4_B5_o , \picorv32_core/sel41_b8/or_B6_B7_o );
  or \picorv32_core/sel41_b8/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [8], \picorv32_core/sel41_b8/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b8/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel41_b9/and_b0_0  (\picorv32_core/sel41_b9/B0 , \picorv32_core/n656 [9], \picorv32_core/n669 );
  and \picorv32_core/sel41_b9/and_b0_1  (\picorv32_core/sel41_b9/B1 , \picorv32_core/n584 [9], \picorv32_core/n668 );
  and \picorv32_core/sel41_b9/and_b0_2  (\picorv32_core/sel41_b9/B2 , \picorv32_core/n570 [9], \picorv32_core/n667 );
  and \picorv32_core/sel41_b9/and_b0_3  (\picorv32_core/sel41_b9/B3 , \picorv32_core/pcpi_rs1$9$ , \picorv32_core/n666 );
  and \picorv32_core/sel41_b9/and_b0_4  (\picorv32_core/sel41_b9/B4 , \picorv32_core/pcpi_rs1$9$ , \picorv32_core/n665 );
  and \picorv32_core/sel41_b9/and_b0_5  (\picorv32_core/sel41_b9/B5 , \picorv32_core/n527 [9], \picorv32_core/n664 );
  and \picorv32_core/sel41_b9/and_b0_6  (\picorv32_core/sel41_b9/B6 , \picorv32_core/pcpi_rs1$9$ , \picorv32_core/n663 );
  and \picorv32_core/sel41_b9/and_b0_7  (\picorv32_core/sel41_b9/B7 , \picorv32_core/pcpi_rs1$9$ , \picorv32_core/n662 );
  or \picorv32_core/sel41_b9/or_B0_B1  (\picorv32_core/sel41_b9/or_B0_B1_o , \picorv32_core/sel41_b9/B0 , \picorv32_core/sel41_b9/B1 );
  or \picorv32_core/sel41_b9/or_B2_B3  (\picorv32_core/sel41_b9/or_B2_B3_o , \picorv32_core/sel41_b9/B2 , \picorv32_core/sel41_b9/B3 );
  or \picorv32_core/sel41_b9/or_B4_B5  (\picorv32_core/sel41_b9/or_B4_B5_o , \picorv32_core/sel41_b9/B4 , \picorv32_core/sel41_b9/B5 );
  or \picorv32_core/sel41_b9/or_B6_B7  (\picorv32_core/sel41_b9/or_B6_B7_o , \picorv32_core/sel41_b9/B6 , \picorv32_core/sel41_b9/B7 );
  or \picorv32_core/sel41_b9/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel41_b9/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b9/or_B0_B1_o , \picorv32_core/sel41_b9/or_B2_B3_o );
  or \picorv32_core/sel41_b9/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel41_b9/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel41_b9/or_B4_B5_o , \picorv32_core/sel41_b9/or_B6_B7_o );
  or \picorv32_core/sel41_b9/or_or_or_B0_B1_o_or_  (\picorv32_core/n693 [9], \picorv32_core/sel41_b9/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel41_b9/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b0/and_b0_0  (\picorv32_core/sel42_b0/B0 , mem_la_wdata[0], \picorv32_core/n669 );
  and \picorv32_core/sel42_b0/and_b0_1  (\picorv32_core/sel42_b0/B1 , mem_la_wdata[0], \picorv32_core/n668 );
  and \picorv32_core/sel42_b0/and_b0_2  (\picorv32_core/sel42_b0/B2 , mem_la_wdata[0], \picorv32_core/n667 );
  and \picorv32_core/sel42_b0/and_b0_3  (\picorv32_core/sel42_b0/B3 , mem_la_wdata[0], \picorv32_core/n666 );
  and \picorv32_core/sel42_b0/and_b0_4  (\picorv32_core/sel42_b0/B4 , \picorv32_core/cpuregs_rs2 [0], \picorv32_core/n665 );
  and \picorv32_core/sel42_b0/and_b0_5  (\picorv32_core/sel42_b0/B5 , \picorv32_core/n528 [0], \picorv32_core/n664 );
  and \picorv32_core/sel42_b0/and_b0_6  (\picorv32_core/sel42_b0/B6 , mem_la_wdata[0], \picorv32_core/n663 );
  and \picorv32_core/sel42_b0/and_b0_7  (\picorv32_core/sel42_b0/B7 , mem_la_wdata[0], \picorv32_core/n662 );
  or \picorv32_core/sel42_b0/or_B0_B1  (\picorv32_core/sel42_b0/or_B0_B1_o , \picorv32_core/sel42_b0/B0 , \picorv32_core/sel42_b0/B1 );
  or \picorv32_core/sel42_b0/or_B2_B3  (\picorv32_core/sel42_b0/or_B2_B3_o , \picorv32_core/sel42_b0/B2 , \picorv32_core/sel42_b0/B3 );
  or \picorv32_core/sel42_b0/or_B4_B5  (\picorv32_core/sel42_b0/or_B4_B5_o , \picorv32_core/sel42_b0/B4 , \picorv32_core/sel42_b0/B5 );
  or \picorv32_core/sel42_b0/or_B6_B7  (\picorv32_core/sel42_b0/or_B6_B7_o , \picorv32_core/sel42_b0/B6 , \picorv32_core/sel42_b0/B7 );
  or \picorv32_core/sel42_b0/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b0/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b0/or_B0_B1_o , \picorv32_core/sel42_b0/or_B2_B3_o );
  or \picorv32_core/sel42_b0/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b0/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b0/or_B4_B5_o , \picorv32_core/sel42_b0/or_B6_B7_o );
  or \picorv32_core/sel42_b0/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [0], \picorv32_core/sel42_b0/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b0/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b1/and_b0_0  (\picorv32_core/sel42_b1/B0 , mem_la_wdata[1], \picorv32_core/n669 );
  and \picorv32_core/sel42_b1/and_b0_1  (\picorv32_core/sel42_b1/B1 , mem_la_wdata[1], \picorv32_core/n668 );
  and \picorv32_core/sel42_b1/and_b0_2  (\picorv32_core/sel42_b1/B2 , mem_la_wdata[1], \picorv32_core/n667 );
  and \picorv32_core/sel42_b1/and_b0_3  (\picorv32_core/sel42_b1/B3 , mem_la_wdata[1], \picorv32_core/n666 );
  and \picorv32_core/sel42_b1/and_b0_4  (\picorv32_core/sel42_b1/B4 , \picorv32_core/cpuregs_rs2 [1], \picorv32_core/n665 );
  and \picorv32_core/sel42_b1/and_b0_5  (\picorv32_core/sel42_b1/B5 , \picorv32_core/n528 [1], \picorv32_core/n664 );
  and \picorv32_core/sel42_b1/and_b0_6  (\picorv32_core/sel42_b1/B6 , mem_la_wdata[1], \picorv32_core/n663 );
  and \picorv32_core/sel42_b1/and_b0_7  (\picorv32_core/sel42_b1/B7 , mem_la_wdata[1], \picorv32_core/n662 );
  or \picorv32_core/sel42_b1/or_B0_B1  (\picorv32_core/sel42_b1/or_B0_B1_o , \picorv32_core/sel42_b1/B0 , \picorv32_core/sel42_b1/B1 );
  or \picorv32_core/sel42_b1/or_B2_B3  (\picorv32_core/sel42_b1/or_B2_B3_o , \picorv32_core/sel42_b1/B2 , \picorv32_core/sel42_b1/B3 );
  or \picorv32_core/sel42_b1/or_B4_B5  (\picorv32_core/sel42_b1/or_B4_B5_o , \picorv32_core/sel42_b1/B4 , \picorv32_core/sel42_b1/B5 );
  or \picorv32_core/sel42_b1/or_B6_B7  (\picorv32_core/sel42_b1/or_B6_B7_o , \picorv32_core/sel42_b1/B6 , \picorv32_core/sel42_b1/B7 );
  or \picorv32_core/sel42_b1/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b1/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b1/or_B0_B1_o , \picorv32_core/sel42_b1/or_B2_B3_o );
  or \picorv32_core/sel42_b1/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b1/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b1/or_B4_B5_o , \picorv32_core/sel42_b1/or_B6_B7_o );
  or \picorv32_core/sel42_b1/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [1], \picorv32_core/sel42_b1/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b1/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b10/and_b0_0  (\picorv32_core/sel42_b10/B0 , \picorv32_core/pcpi_rs2$10$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b10/and_b0_1  (\picorv32_core/sel42_b10/B1 , \picorv32_core/pcpi_rs2$10$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b10/and_b0_2  (\picorv32_core/sel42_b10/B2 , \picorv32_core/pcpi_rs2$10$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b10/and_b0_3  (\picorv32_core/sel42_b10/B3 , \picorv32_core/pcpi_rs2$10$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b10/and_b0_4  (\picorv32_core/sel42_b10/B4 , \picorv32_core/cpuregs_rs2 [10], \picorv32_core/n665 );
  and \picorv32_core/sel42_b10/and_b0_5  (\picorv32_core/sel42_b10/B5 , \picorv32_core/n528 [10], \picorv32_core/n664 );
  and \picorv32_core/sel42_b10/and_b0_6  (\picorv32_core/sel42_b10/B6 , \picorv32_core/pcpi_rs2$10$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b10/and_b0_7  (\picorv32_core/sel42_b10/B7 , \picorv32_core/pcpi_rs2$10$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b10/or_B0_B1  (\picorv32_core/sel42_b10/or_B0_B1_o , \picorv32_core/sel42_b10/B0 , \picorv32_core/sel42_b10/B1 );
  or \picorv32_core/sel42_b10/or_B2_B3  (\picorv32_core/sel42_b10/or_B2_B3_o , \picorv32_core/sel42_b10/B2 , \picorv32_core/sel42_b10/B3 );
  or \picorv32_core/sel42_b10/or_B4_B5  (\picorv32_core/sel42_b10/or_B4_B5_o , \picorv32_core/sel42_b10/B4 , \picorv32_core/sel42_b10/B5 );
  or \picorv32_core/sel42_b10/or_B6_B7  (\picorv32_core/sel42_b10/or_B6_B7_o , \picorv32_core/sel42_b10/B6 , \picorv32_core/sel42_b10/B7 );
  or \picorv32_core/sel42_b10/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b10/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b10/or_B0_B1_o , \picorv32_core/sel42_b10/or_B2_B3_o );
  or \picorv32_core/sel42_b10/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b10/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b10/or_B4_B5_o , \picorv32_core/sel42_b10/or_B6_B7_o );
  or \picorv32_core/sel42_b10/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [10], \picorv32_core/sel42_b10/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b10/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b11/and_b0_0  (\picorv32_core/sel42_b11/B0 , \picorv32_core/pcpi_rs2$11$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b11/and_b0_1  (\picorv32_core/sel42_b11/B1 , \picorv32_core/pcpi_rs2$11$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b11/and_b0_2  (\picorv32_core/sel42_b11/B2 , \picorv32_core/pcpi_rs2$11$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b11/and_b0_3  (\picorv32_core/sel42_b11/B3 , \picorv32_core/pcpi_rs2$11$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b11/and_b0_4  (\picorv32_core/sel42_b11/B4 , \picorv32_core/cpuregs_rs2 [11], \picorv32_core/n665 );
  and \picorv32_core/sel42_b11/and_b0_5  (\picorv32_core/sel42_b11/B5 , \picorv32_core/n528 [11], \picorv32_core/n664 );
  and \picorv32_core/sel42_b11/and_b0_6  (\picorv32_core/sel42_b11/B6 , \picorv32_core/pcpi_rs2$11$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b11/and_b0_7  (\picorv32_core/sel42_b11/B7 , \picorv32_core/pcpi_rs2$11$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b11/or_B0_B1  (\picorv32_core/sel42_b11/or_B0_B1_o , \picorv32_core/sel42_b11/B0 , \picorv32_core/sel42_b11/B1 );
  or \picorv32_core/sel42_b11/or_B2_B3  (\picorv32_core/sel42_b11/or_B2_B3_o , \picorv32_core/sel42_b11/B2 , \picorv32_core/sel42_b11/B3 );
  or \picorv32_core/sel42_b11/or_B4_B5  (\picorv32_core/sel42_b11/or_B4_B5_o , \picorv32_core/sel42_b11/B4 , \picorv32_core/sel42_b11/B5 );
  or \picorv32_core/sel42_b11/or_B6_B7  (\picorv32_core/sel42_b11/or_B6_B7_o , \picorv32_core/sel42_b11/B6 , \picorv32_core/sel42_b11/B7 );
  or \picorv32_core/sel42_b11/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b11/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b11/or_B0_B1_o , \picorv32_core/sel42_b11/or_B2_B3_o );
  or \picorv32_core/sel42_b11/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b11/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b11/or_B4_B5_o , \picorv32_core/sel42_b11/or_B6_B7_o );
  or \picorv32_core/sel42_b11/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [11], \picorv32_core/sel42_b11/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b11/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b12/and_b0_0  (\picorv32_core/sel42_b12/B0 , \picorv32_core/pcpi_rs2$12$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b12/and_b0_1  (\picorv32_core/sel42_b12/B1 , \picorv32_core/pcpi_rs2$12$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b12/and_b0_2  (\picorv32_core/sel42_b12/B2 , \picorv32_core/pcpi_rs2$12$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b12/and_b0_3  (\picorv32_core/sel42_b12/B3 , \picorv32_core/pcpi_rs2$12$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b12/and_b0_4  (\picorv32_core/sel42_b12/B4 , \picorv32_core/cpuregs_rs2 [12], \picorv32_core/n665 );
  and \picorv32_core/sel42_b12/and_b0_5  (\picorv32_core/sel42_b12/B5 , \picorv32_core/n528 [12], \picorv32_core/n664 );
  and \picorv32_core/sel42_b12/and_b0_6  (\picorv32_core/sel42_b12/B6 , \picorv32_core/pcpi_rs2$12$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b12/and_b0_7  (\picorv32_core/sel42_b12/B7 , \picorv32_core/pcpi_rs2$12$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b12/or_B0_B1  (\picorv32_core/sel42_b12/or_B0_B1_o , \picorv32_core/sel42_b12/B0 , \picorv32_core/sel42_b12/B1 );
  or \picorv32_core/sel42_b12/or_B2_B3  (\picorv32_core/sel42_b12/or_B2_B3_o , \picorv32_core/sel42_b12/B2 , \picorv32_core/sel42_b12/B3 );
  or \picorv32_core/sel42_b12/or_B4_B5  (\picorv32_core/sel42_b12/or_B4_B5_o , \picorv32_core/sel42_b12/B4 , \picorv32_core/sel42_b12/B5 );
  or \picorv32_core/sel42_b12/or_B6_B7  (\picorv32_core/sel42_b12/or_B6_B7_o , \picorv32_core/sel42_b12/B6 , \picorv32_core/sel42_b12/B7 );
  or \picorv32_core/sel42_b12/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b12/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b12/or_B0_B1_o , \picorv32_core/sel42_b12/or_B2_B3_o );
  or \picorv32_core/sel42_b12/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b12/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b12/or_B4_B5_o , \picorv32_core/sel42_b12/or_B6_B7_o );
  or \picorv32_core/sel42_b12/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [12], \picorv32_core/sel42_b12/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b12/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b13/and_b0_0  (\picorv32_core/sel42_b13/B0 , \picorv32_core/pcpi_rs2$13$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b13/and_b0_1  (\picorv32_core/sel42_b13/B1 , \picorv32_core/pcpi_rs2$13$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b13/and_b0_2  (\picorv32_core/sel42_b13/B2 , \picorv32_core/pcpi_rs2$13$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b13/and_b0_3  (\picorv32_core/sel42_b13/B3 , \picorv32_core/pcpi_rs2$13$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b13/and_b0_4  (\picorv32_core/sel42_b13/B4 , \picorv32_core/cpuregs_rs2 [13], \picorv32_core/n665 );
  and \picorv32_core/sel42_b13/and_b0_5  (\picorv32_core/sel42_b13/B5 , \picorv32_core/n528 [13], \picorv32_core/n664 );
  and \picorv32_core/sel42_b13/and_b0_6  (\picorv32_core/sel42_b13/B6 , \picorv32_core/pcpi_rs2$13$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b13/and_b0_7  (\picorv32_core/sel42_b13/B7 , \picorv32_core/pcpi_rs2$13$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b13/or_B0_B1  (\picorv32_core/sel42_b13/or_B0_B1_o , \picorv32_core/sel42_b13/B0 , \picorv32_core/sel42_b13/B1 );
  or \picorv32_core/sel42_b13/or_B2_B3  (\picorv32_core/sel42_b13/or_B2_B3_o , \picorv32_core/sel42_b13/B2 , \picorv32_core/sel42_b13/B3 );
  or \picorv32_core/sel42_b13/or_B4_B5  (\picorv32_core/sel42_b13/or_B4_B5_o , \picorv32_core/sel42_b13/B4 , \picorv32_core/sel42_b13/B5 );
  or \picorv32_core/sel42_b13/or_B6_B7  (\picorv32_core/sel42_b13/or_B6_B7_o , \picorv32_core/sel42_b13/B6 , \picorv32_core/sel42_b13/B7 );
  or \picorv32_core/sel42_b13/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b13/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b13/or_B0_B1_o , \picorv32_core/sel42_b13/or_B2_B3_o );
  or \picorv32_core/sel42_b13/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b13/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b13/or_B4_B5_o , \picorv32_core/sel42_b13/or_B6_B7_o );
  or \picorv32_core/sel42_b13/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [13], \picorv32_core/sel42_b13/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b13/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b14/and_b0_0  (\picorv32_core/sel42_b14/B0 , \picorv32_core/pcpi_rs2$14$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b14/and_b0_1  (\picorv32_core/sel42_b14/B1 , \picorv32_core/pcpi_rs2$14$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b14/and_b0_2  (\picorv32_core/sel42_b14/B2 , \picorv32_core/pcpi_rs2$14$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b14/and_b0_3  (\picorv32_core/sel42_b14/B3 , \picorv32_core/pcpi_rs2$14$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b14/and_b0_4  (\picorv32_core/sel42_b14/B4 , \picorv32_core/cpuregs_rs2 [14], \picorv32_core/n665 );
  and \picorv32_core/sel42_b14/and_b0_5  (\picorv32_core/sel42_b14/B5 , \picorv32_core/n528 [14], \picorv32_core/n664 );
  and \picorv32_core/sel42_b14/and_b0_6  (\picorv32_core/sel42_b14/B6 , \picorv32_core/pcpi_rs2$14$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b14/and_b0_7  (\picorv32_core/sel42_b14/B7 , \picorv32_core/pcpi_rs2$14$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b14/or_B0_B1  (\picorv32_core/sel42_b14/or_B0_B1_o , \picorv32_core/sel42_b14/B0 , \picorv32_core/sel42_b14/B1 );
  or \picorv32_core/sel42_b14/or_B2_B3  (\picorv32_core/sel42_b14/or_B2_B3_o , \picorv32_core/sel42_b14/B2 , \picorv32_core/sel42_b14/B3 );
  or \picorv32_core/sel42_b14/or_B4_B5  (\picorv32_core/sel42_b14/or_B4_B5_o , \picorv32_core/sel42_b14/B4 , \picorv32_core/sel42_b14/B5 );
  or \picorv32_core/sel42_b14/or_B6_B7  (\picorv32_core/sel42_b14/or_B6_B7_o , \picorv32_core/sel42_b14/B6 , \picorv32_core/sel42_b14/B7 );
  or \picorv32_core/sel42_b14/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b14/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b14/or_B0_B1_o , \picorv32_core/sel42_b14/or_B2_B3_o );
  or \picorv32_core/sel42_b14/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b14/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b14/or_B4_B5_o , \picorv32_core/sel42_b14/or_B6_B7_o );
  or \picorv32_core/sel42_b14/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [14], \picorv32_core/sel42_b14/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b14/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b15/and_b0_0  (\picorv32_core/sel42_b15/B0 , \picorv32_core/pcpi_rs2$15$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b15/and_b0_1  (\picorv32_core/sel42_b15/B1 , \picorv32_core/pcpi_rs2$15$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b15/and_b0_2  (\picorv32_core/sel42_b15/B2 , \picorv32_core/pcpi_rs2$15$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b15/and_b0_3  (\picorv32_core/sel42_b15/B3 , \picorv32_core/pcpi_rs2$15$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b15/and_b0_4  (\picorv32_core/sel42_b15/B4 , \picorv32_core/cpuregs_rs2 [15], \picorv32_core/n665 );
  and \picorv32_core/sel42_b15/and_b0_5  (\picorv32_core/sel42_b15/B5 , \picorv32_core/n528 [15], \picorv32_core/n664 );
  and \picorv32_core/sel42_b15/and_b0_6  (\picorv32_core/sel42_b15/B6 , \picorv32_core/pcpi_rs2$15$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b15/and_b0_7  (\picorv32_core/sel42_b15/B7 , \picorv32_core/pcpi_rs2$15$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b15/or_B0_B1  (\picorv32_core/sel42_b15/or_B0_B1_o , \picorv32_core/sel42_b15/B0 , \picorv32_core/sel42_b15/B1 );
  or \picorv32_core/sel42_b15/or_B2_B3  (\picorv32_core/sel42_b15/or_B2_B3_o , \picorv32_core/sel42_b15/B2 , \picorv32_core/sel42_b15/B3 );
  or \picorv32_core/sel42_b15/or_B4_B5  (\picorv32_core/sel42_b15/or_B4_B5_o , \picorv32_core/sel42_b15/B4 , \picorv32_core/sel42_b15/B5 );
  or \picorv32_core/sel42_b15/or_B6_B7  (\picorv32_core/sel42_b15/or_B6_B7_o , \picorv32_core/sel42_b15/B6 , \picorv32_core/sel42_b15/B7 );
  or \picorv32_core/sel42_b15/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b15/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b15/or_B0_B1_o , \picorv32_core/sel42_b15/or_B2_B3_o );
  or \picorv32_core/sel42_b15/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b15/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b15/or_B4_B5_o , \picorv32_core/sel42_b15/or_B6_B7_o );
  or \picorv32_core/sel42_b15/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [15], \picorv32_core/sel42_b15/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b15/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b16/and_b0_0  (\picorv32_core/sel42_b16/B0 , \picorv32_core/pcpi_rs2$16$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b16/and_b0_1  (\picorv32_core/sel42_b16/B1 , \picorv32_core/pcpi_rs2$16$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b16/and_b0_2  (\picorv32_core/sel42_b16/B2 , \picorv32_core/pcpi_rs2$16$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b16/and_b0_3  (\picorv32_core/sel42_b16/B3 , \picorv32_core/pcpi_rs2$16$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b16/and_b0_4  (\picorv32_core/sel42_b16/B4 , \picorv32_core/cpuregs_rs2 [16], \picorv32_core/n665 );
  and \picorv32_core/sel42_b16/and_b0_5  (\picorv32_core/sel42_b16/B5 , \picorv32_core/n528 [16], \picorv32_core/n664 );
  and \picorv32_core/sel42_b16/and_b0_6  (\picorv32_core/sel42_b16/B6 , \picorv32_core/pcpi_rs2$16$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b16/and_b0_7  (\picorv32_core/sel42_b16/B7 , \picorv32_core/pcpi_rs2$16$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b16/or_B0_B1  (\picorv32_core/sel42_b16/or_B0_B1_o , \picorv32_core/sel42_b16/B0 , \picorv32_core/sel42_b16/B1 );
  or \picorv32_core/sel42_b16/or_B2_B3  (\picorv32_core/sel42_b16/or_B2_B3_o , \picorv32_core/sel42_b16/B2 , \picorv32_core/sel42_b16/B3 );
  or \picorv32_core/sel42_b16/or_B4_B5  (\picorv32_core/sel42_b16/or_B4_B5_o , \picorv32_core/sel42_b16/B4 , \picorv32_core/sel42_b16/B5 );
  or \picorv32_core/sel42_b16/or_B6_B7  (\picorv32_core/sel42_b16/or_B6_B7_o , \picorv32_core/sel42_b16/B6 , \picorv32_core/sel42_b16/B7 );
  or \picorv32_core/sel42_b16/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b16/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b16/or_B0_B1_o , \picorv32_core/sel42_b16/or_B2_B3_o );
  or \picorv32_core/sel42_b16/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b16/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b16/or_B4_B5_o , \picorv32_core/sel42_b16/or_B6_B7_o );
  or \picorv32_core/sel42_b16/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [16], \picorv32_core/sel42_b16/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b16/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b17/and_b0_0  (\picorv32_core/sel42_b17/B0 , \picorv32_core/pcpi_rs2$17$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b17/and_b0_1  (\picorv32_core/sel42_b17/B1 , \picorv32_core/pcpi_rs2$17$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b17/and_b0_2  (\picorv32_core/sel42_b17/B2 , \picorv32_core/pcpi_rs2$17$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b17/and_b0_3  (\picorv32_core/sel42_b17/B3 , \picorv32_core/pcpi_rs2$17$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b17/and_b0_4  (\picorv32_core/sel42_b17/B4 , \picorv32_core/cpuregs_rs2 [17], \picorv32_core/n665 );
  and \picorv32_core/sel42_b17/and_b0_5  (\picorv32_core/sel42_b17/B5 , \picorv32_core/n528 [17], \picorv32_core/n664 );
  and \picorv32_core/sel42_b17/and_b0_6  (\picorv32_core/sel42_b17/B6 , \picorv32_core/pcpi_rs2$17$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b17/and_b0_7  (\picorv32_core/sel42_b17/B7 , \picorv32_core/pcpi_rs2$17$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b17/or_B0_B1  (\picorv32_core/sel42_b17/or_B0_B1_o , \picorv32_core/sel42_b17/B0 , \picorv32_core/sel42_b17/B1 );
  or \picorv32_core/sel42_b17/or_B2_B3  (\picorv32_core/sel42_b17/or_B2_B3_o , \picorv32_core/sel42_b17/B2 , \picorv32_core/sel42_b17/B3 );
  or \picorv32_core/sel42_b17/or_B4_B5  (\picorv32_core/sel42_b17/or_B4_B5_o , \picorv32_core/sel42_b17/B4 , \picorv32_core/sel42_b17/B5 );
  or \picorv32_core/sel42_b17/or_B6_B7  (\picorv32_core/sel42_b17/or_B6_B7_o , \picorv32_core/sel42_b17/B6 , \picorv32_core/sel42_b17/B7 );
  or \picorv32_core/sel42_b17/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b17/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b17/or_B0_B1_o , \picorv32_core/sel42_b17/or_B2_B3_o );
  or \picorv32_core/sel42_b17/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b17/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b17/or_B4_B5_o , \picorv32_core/sel42_b17/or_B6_B7_o );
  or \picorv32_core/sel42_b17/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [17], \picorv32_core/sel42_b17/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b17/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b18/and_b0_0  (\picorv32_core/sel42_b18/B0 , \picorv32_core/pcpi_rs2$18$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b18/and_b0_1  (\picorv32_core/sel42_b18/B1 , \picorv32_core/pcpi_rs2$18$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b18/and_b0_2  (\picorv32_core/sel42_b18/B2 , \picorv32_core/pcpi_rs2$18$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b18/and_b0_3  (\picorv32_core/sel42_b18/B3 , \picorv32_core/pcpi_rs2$18$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b18/and_b0_4  (\picorv32_core/sel42_b18/B4 , \picorv32_core/cpuregs_rs2 [18], \picorv32_core/n665 );
  and \picorv32_core/sel42_b18/and_b0_5  (\picorv32_core/sel42_b18/B5 , \picorv32_core/n528 [18], \picorv32_core/n664 );
  and \picorv32_core/sel42_b18/and_b0_6  (\picorv32_core/sel42_b18/B6 , \picorv32_core/pcpi_rs2$18$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b18/and_b0_7  (\picorv32_core/sel42_b18/B7 , \picorv32_core/pcpi_rs2$18$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b18/or_B0_B1  (\picorv32_core/sel42_b18/or_B0_B1_o , \picorv32_core/sel42_b18/B0 , \picorv32_core/sel42_b18/B1 );
  or \picorv32_core/sel42_b18/or_B2_B3  (\picorv32_core/sel42_b18/or_B2_B3_o , \picorv32_core/sel42_b18/B2 , \picorv32_core/sel42_b18/B3 );
  or \picorv32_core/sel42_b18/or_B4_B5  (\picorv32_core/sel42_b18/or_B4_B5_o , \picorv32_core/sel42_b18/B4 , \picorv32_core/sel42_b18/B5 );
  or \picorv32_core/sel42_b18/or_B6_B7  (\picorv32_core/sel42_b18/or_B6_B7_o , \picorv32_core/sel42_b18/B6 , \picorv32_core/sel42_b18/B7 );
  or \picorv32_core/sel42_b18/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b18/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b18/or_B0_B1_o , \picorv32_core/sel42_b18/or_B2_B3_o );
  or \picorv32_core/sel42_b18/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b18/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b18/or_B4_B5_o , \picorv32_core/sel42_b18/or_B6_B7_o );
  or \picorv32_core/sel42_b18/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [18], \picorv32_core/sel42_b18/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b18/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b19/and_b0_0  (\picorv32_core/sel42_b19/B0 , \picorv32_core/pcpi_rs2$19$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b19/and_b0_1  (\picorv32_core/sel42_b19/B1 , \picorv32_core/pcpi_rs2$19$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b19/and_b0_2  (\picorv32_core/sel42_b19/B2 , \picorv32_core/pcpi_rs2$19$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b19/and_b0_3  (\picorv32_core/sel42_b19/B3 , \picorv32_core/pcpi_rs2$19$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b19/and_b0_4  (\picorv32_core/sel42_b19/B4 , \picorv32_core/cpuregs_rs2 [19], \picorv32_core/n665 );
  and \picorv32_core/sel42_b19/and_b0_5  (\picorv32_core/sel42_b19/B5 , \picorv32_core/n528 [19], \picorv32_core/n664 );
  and \picorv32_core/sel42_b19/and_b0_6  (\picorv32_core/sel42_b19/B6 , \picorv32_core/pcpi_rs2$19$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b19/and_b0_7  (\picorv32_core/sel42_b19/B7 , \picorv32_core/pcpi_rs2$19$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b19/or_B0_B1  (\picorv32_core/sel42_b19/or_B0_B1_o , \picorv32_core/sel42_b19/B0 , \picorv32_core/sel42_b19/B1 );
  or \picorv32_core/sel42_b19/or_B2_B3  (\picorv32_core/sel42_b19/or_B2_B3_o , \picorv32_core/sel42_b19/B2 , \picorv32_core/sel42_b19/B3 );
  or \picorv32_core/sel42_b19/or_B4_B5  (\picorv32_core/sel42_b19/or_B4_B5_o , \picorv32_core/sel42_b19/B4 , \picorv32_core/sel42_b19/B5 );
  or \picorv32_core/sel42_b19/or_B6_B7  (\picorv32_core/sel42_b19/or_B6_B7_o , \picorv32_core/sel42_b19/B6 , \picorv32_core/sel42_b19/B7 );
  or \picorv32_core/sel42_b19/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b19/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b19/or_B0_B1_o , \picorv32_core/sel42_b19/or_B2_B3_o );
  or \picorv32_core/sel42_b19/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b19/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b19/or_B4_B5_o , \picorv32_core/sel42_b19/or_B6_B7_o );
  or \picorv32_core/sel42_b19/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [19], \picorv32_core/sel42_b19/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b19/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b2/and_b0_0  (\picorv32_core/sel42_b2/B0 , mem_la_wdata[2], \picorv32_core/n669 );
  and \picorv32_core/sel42_b2/and_b0_1  (\picorv32_core/sel42_b2/B1 , mem_la_wdata[2], \picorv32_core/n668 );
  and \picorv32_core/sel42_b2/and_b0_2  (\picorv32_core/sel42_b2/B2 , mem_la_wdata[2], \picorv32_core/n667 );
  and \picorv32_core/sel42_b2/and_b0_3  (\picorv32_core/sel42_b2/B3 , mem_la_wdata[2], \picorv32_core/n666 );
  and \picorv32_core/sel42_b2/and_b0_4  (\picorv32_core/sel42_b2/B4 , \picorv32_core/cpuregs_rs2 [2], \picorv32_core/n665 );
  and \picorv32_core/sel42_b2/and_b0_5  (\picorv32_core/sel42_b2/B5 , \picorv32_core/n528 [2], \picorv32_core/n664 );
  and \picorv32_core/sel42_b2/and_b0_6  (\picorv32_core/sel42_b2/B6 , mem_la_wdata[2], \picorv32_core/n663 );
  and \picorv32_core/sel42_b2/and_b0_7  (\picorv32_core/sel42_b2/B7 , mem_la_wdata[2], \picorv32_core/n662 );
  or \picorv32_core/sel42_b2/or_B0_B1  (\picorv32_core/sel42_b2/or_B0_B1_o , \picorv32_core/sel42_b2/B0 , \picorv32_core/sel42_b2/B1 );
  or \picorv32_core/sel42_b2/or_B2_B3  (\picorv32_core/sel42_b2/or_B2_B3_o , \picorv32_core/sel42_b2/B2 , \picorv32_core/sel42_b2/B3 );
  or \picorv32_core/sel42_b2/or_B4_B5  (\picorv32_core/sel42_b2/or_B4_B5_o , \picorv32_core/sel42_b2/B4 , \picorv32_core/sel42_b2/B5 );
  or \picorv32_core/sel42_b2/or_B6_B7  (\picorv32_core/sel42_b2/or_B6_B7_o , \picorv32_core/sel42_b2/B6 , \picorv32_core/sel42_b2/B7 );
  or \picorv32_core/sel42_b2/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b2/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b2/or_B0_B1_o , \picorv32_core/sel42_b2/or_B2_B3_o );
  or \picorv32_core/sel42_b2/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b2/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b2/or_B4_B5_o , \picorv32_core/sel42_b2/or_B6_B7_o );
  or \picorv32_core/sel42_b2/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [2], \picorv32_core/sel42_b2/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b2/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b20/and_b0_0  (\picorv32_core/sel42_b20/B0 , \picorv32_core/pcpi_rs2$20$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b20/and_b0_1  (\picorv32_core/sel42_b20/B1 , \picorv32_core/pcpi_rs2$20$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b20/and_b0_2  (\picorv32_core/sel42_b20/B2 , \picorv32_core/pcpi_rs2$20$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b20/and_b0_3  (\picorv32_core/sel42_b20/B3 , \picorv32_core/pcpi_rs2$20$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b20/and_b0_4  (\picorv32_core/sel42_b20/B4 , \picorv32_core/cpuregs_rs2 [20], \picorv32_core/n665 );
  and \picorv32_core/sel42_b20/and_b0_5  (\picorv32_core/sel42_b20/B5 , \picorv32_core/n528 [20], \picorv32_core/n664 );
  and \picorv32_core/sel42_b20/and_b0_6  (\picorv32_core/sel42_b20/B6 , \picorv32_core/pcpi_rs2$20$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b20/and_b0_7  (\picorv32_core/sel42_b20/B7 , \picorv32_core/pcpi_rs2$20$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b20/or_B0_B1  (\picorv32_core/sel42_b20/or_B0_B1_o , \picorv32_core/sel42_b20/B0 , \picorv32_core/sel42_b20/B1 );
  or \picorv32_core/sel42_b20/or_B2_B3  (\picorv32_core/sel42_b20/or_B2_B3_o , \picorv32_core/sel42_b20/B2 , \picorv32_core/sel42_b20/B3 );
  or \picorv32_core/sel42_b20/or_B4_B5  (\picorv32_core/sel42_b20/or_B4_B5_o , \picorv32_core/sel42_b20/B4 , \picorv32_core/sel42_b20/B5 );
  or \picorv32_core/sel42_b20/or_B6_B7  (\picorv32_core/sel42_b20/or_B6_B7_o , \picorv32_core/sel42_b20/B6 , \picorv32_core/sel42_b20/B7 );
  or \picorv32_core/sel42_b20/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b20/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b20/or_B0_B1_o , \picorv32_core/sel42_b20/or_B2_B3_o );
  or \picorv32_core/sel42_b20/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b20/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b20/or_B4_B5_o , \picorv32_core/sel42_b20/or_B6_B7_o );
  or \picorv32_core/sel42_b20/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [20], \picorv32_core/sel42_b20/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b20/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b21/and_b0_0  (\picorv32_core/sel42_b21/B0 , \picorv32_core/pcpi_rs2$21$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b21/and_b0_1  (\picorv32_core/sel42_b21/B1 , \picorv32_core/pcpi_rs2$21$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b21/and_b0_2  (\picorv32_core/sel42_b21/B2 , \picorv32_core/pcpi_rs2$21$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b21/and_b0_3  (\picorv32_core/sel42_b21/B3 , \picorv32_core/pcpi_rs2$21$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b21/and_b0_4  (\picorv32_core/sel42_b21/B4 , \picorv32_core/cpuregs_rs2 [21], \picorv32_core/n665 );
  and \picorv32_core/sel42_b21/and_b0_5  (\picorv32_core/sel42_b21/B5 , \picorv32_core/n528 [21], \picorv32_core/n664 );
  and \picorv32_core/sel42_b21/and_b0_6  (\picorv32_core/sel42_b21/B6 , \picorv32_core/pcpi_rs2$21$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b21/and_b0_7  (\picorv32_core/sel42_b21/B7 , \picorv32_core/pcpi_rs2$21$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b21/or_B0_B1  (\picorv32_core/sel42_b21/or_B0_B1_o , \picorv32_core/sel42_b21/B0 , \picorv32_core/sel42_b21/B1 );
  or \picorv32_core/sel42_b21/or_B2_B3  (\picorv32_core/sel42_b21/or_B2_B3_o , \picorv32_core/sel42_b21/B2 , \picorv32_core/sel42_b21/B3 );
  or \picorv32_core/sel42_b21/or_B4_B5  (\picorv32_core/sel42_b21/or_B4_B5_o , \picorv32_core/sel42_b21/B4 , \picorv32_core/sel42_b21/B5 );
  or \picorv32_core/sel42_b21/or_B6_B7  (\picorv32_core/sel42_b21/or_B6_B7_o , \picorv32_core/sel42_b21/B6 , \picorv32_core/sel42_b21/B7 );
  or \picorv32_core/sel42_b21/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b21/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b21/or_B0_B1_o , \picorv32_core/sel42_b21/or_B2_B3_o );
  or \picorv32_core/sel42_b21/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b21/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b21/or_B4_B5_o , \picorv32_core/sel42_b21/or_B6_B7_o );
  or \picorv32_core/sel42_b21/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [21], \picorv32_core/sel42_b21/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b21/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b22/and_b0_0  (\picorv32_core/sel42_b22/B0 , \picorv32_core/pcpi_rs2$22$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b22/and_b0_1  (\picorv32_core/sel42_b22/B1 , \picorv32_core/pcpi_rs2$22$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b22/and_b0_2  (\picorv32_core/sel42_b22/B2 , \picorv32_core/pcpi_rs2$22$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b22/and_b0_3  (\picorv32_core/sel42_b22/B3 , \picorv32_core/pcpi_rs2$22$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b22/and_b0_4  (\picorv32_core/sel42_b22/B4 , \picorv32_core/cpuregs_rs2 [22], \picorv32_core/n665 );
  and \picorv32_core/sel42_b22/and_b0_5  (\picorv32_core/sel42_b22/B5 , \picorv32_core/n528 [22], \picorv32_core/n664 );
  and \picorv32_core/sel42_b22/and_b0_6  (\picorv32_core/sel42_b22/B6 , \picorv32_core/pcpi_rs2$22$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b22/and_b0_7  (\picorv32_core/sel42_b22/B7 , \picorv32_core/pcpi_rs2$22$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b22/or_B0_B1  (\picorv32_core/sel42_b22/or_B0_B1_o , \picorv32_core/sel42_b22/B0 , \picorv32_core/sel42_b22/B1 );
  or \picorv32_core/sel42_b22/or_B2_B3  (\picorv32_core/sel42_b22/or_B2_B3_o , \picorv32_core/sel42_b22/B2 , \picorv32_core/sel42_b22/B3 );
  or \picorv32_core/sel42_b22/or_B4_B5  (\picorv32_core/sel42_b22/or_B4_B5_o , \picorv32_core/sel42_b22/B4 , \picorv32_core/sel42_b22/B5 );
  or \picorv32_core/sel42_b22/or_B6_B7  (\picorv32_core/sel42_b22/or_B6_B7_o , \picorv32_core/sel42_b22/B6 , \picorv32_core/sel42_b22/B7 );
  or \picorv32_core/sel42_b22/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b22/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b22/or_B0_B1_o , \picorv32_core/sel42_b22/or_B2_B3_o );
  or \picorv32_core/sel42_b22/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b22/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b22/or_B4_B5_o , \picorv32_core/sel42_b22/or_B6_B7_o );
  or \picorv32_core/sel42_b22/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [22], \picorv32_core/sel42_b22/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b22/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b23/and_b0_0  (\picorv32_core/sel42_b23/B0 , \picorv32_core/pcpi_rs2$23$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b23/and_b0_1  (\picorv32_core/sel42_b23/B1 , \picorv32_core/pcpi_rs2$23$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b23/and_b0_2  (\picorv32_core/sel42_b23/B2 , \picorv32_core/pcpi_rs2$23$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b23/and_b0_3  (\picorv32_core/sel42_b23/B3 , \picorv32_core/pcpi_rs2$23$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b23/and_b0_4  (\picorv32_core/sel42_b23/B4 , \picorv32_core/cpuregs_rs2 [23], \picorv32_core/n665 );
  and \picorv32_core/sel42_b23/and_b0_5  (\picorv32_core/sel42_b23/B5 , \picorv32_core/n528 [23], \picorv32_core/n664 );
  and \picorv32_core/sel42_b23/and_b0_6  (\picorv32_core/sel42_b23/B6 , \picorv32_core/pcpi_rs2$23$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b23/and_b0_7  (\picorv32_core/sel42_b23/B7 , \picorv32_core/pcpi_rs2$23$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b23/or_B0_B1  (\picorv32_core/sel42_b23/or_B0_B1_o , \picorv32_core/sel42_b23/B0 , \picorv32_core/sel42_b23/B1 );
  or \picorv32_core/sel42_b23/or_B2_B3  (\picorv32_core/sel42_b23/or_B2_B3_o , \picorv32_core/sel42_b23/B2 , \picorv32_core/sel42_b23/B3 );
  or \picorv32_core/sel42_b23/or_B4_B5  (\picorv32_core/sel42_b23/or_B4_B5_o , \picorv32_core/sel42_b23/B4 , \picorv32_core/sel42_b23/B5 );
  or \picorv32_core/sel42_b23/or_B6_B7  (\picorv32_core/sel42_b23/or_B6_B7_o , \picorv32_core/sel42_b23/B6 , \picorv32_core/sel42_b23/B7 );
  or \picorv32_core/sel42_b23/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b23/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b23/or_B0_B1_o , \picorv32_core/sel42_b23/or_B2_B3_o );
  or \picorv32_core/sel42_b23/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b23/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b23/or_B4_B5_o , \picorv32_core/sel42_b23/or_B6_B7_o );
  or \picorv32_core/sel42_b23/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [23], \picorv32_core/sel42_b23/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b23/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b24/and_b0_0  (\picorv32_core/sel42_b24/B0 , \picorv32_core/pcpi_rs2$24$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b24/and_b0_1  (\picorv32_core/sel42_b24/B1 , \picorv32_core/pcpi_rs2$24$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b24/and_b0_2  (\picorv32_core/sel42_b24/B2 , \picorv32_core/pcpi_rs2$24$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b24/and_b0_3  (\picorv32_core/sel42_b24/B3 , \picorv32_core/pcpi_rs2$24$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b24/and_b0_4  (\picorv32_core/sel42_b24/B4 , \picorv32_core/cpuregs_rs2 [24], \picorv32_core/n665 );
  and \picorv32_core/sel42_b24/and_b0_5  (\picorv32_core/sel42_b24/B5 , \picorv32_core/n528 [24], \picorv32_core/n664 );
  and \picorv32_core/sel42_b24/and_b0_6  (\picorv32_core/sel42_b24/B6 , \picorv32_core/pcpi_rs2$24$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b24/and_b0_7  (\picorv32_core/sel42_b24/B7 , \picorv32_core/pcpi_rs2$24$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b24/or_B0_B1  (\picorv32_core/sel42_b24/or_B0_B1_o , \picorv32_core/sel42_b24/B0 , \picorv32_core/sel42_b24/B1 );
  or \picorv32_core/sel42_b24/or_B2_B3  (\picorv32_core/sel42_b24/or_B2_B3_o , \picorv32_core/sel42_b24/B2 , \picorv32_core/sel42_b24/B3 );
  or \picorv32_core/sel42_b24/or_B4_B5  (\picorv32_core/sel42_b24/or_B4_B5_o , \picorv32_core/sel42_b24/B4 , \picorv32_core/sel42_b24/B5 );
  or \picorv32_core/sel42_b24/or_B6_B7  (\picorv32_core/sel42_b24/or_B6_B7_o , \picorv32_core/sel42_b24/B6 , \picorv32_core/sel42_b24/B7 );
  or \picorv32_core/sel42_b24/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b24/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b24/or_B0_B1_o , \picorv32_core/sel42_b24/or_B2_B3_o );
  or \picorv32_core/sel42_b24/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b24/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b24/or_B4_B5_o , \picorv32_core/sel42_b24/or_B6_B7_o );
  or \picorv32_core/sel42_b24/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [24], \picorv32_core/sel42_b24/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b24/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b25/and_b0_0  (\picorv32_core/sel42_b25/B0 , \picorv32_core/pcpi_rs2$25$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b25/and_b0_1  (\picorv32_core/sel42_b25/B1 , \picorv32_core/pcpi_rs2$25$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b25/and_b0_2  (\picorv32_core/sel42_b25/B2 , \picorv32_core/pcpi_rs2$25$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b25/and_b0_3  (\picorv32_core/sel42_b25/B3 , \picorv32_core/pcpi_rs2$25$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b25/and_b0_4  (\picorv32_core/sel42_b25/B4 , \picorv32_core/cpuregs_rs2 [25], \picorv32_core/n665 );
  and \picorv32_core/sel42_b25/and_b0_5  (\picorv32_core/sel42_b25/B5 , \picorv32_core/n528 [25], \picorv32_core/n664 );
  and \picorv32_core/sel42_b25/and_b0_6  (\picorv32_core/sel42_b25/B6 , \picorv32_core/pcpi_rs2$25$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b25/and_b0_7  (\picorv32_core/sel42_b25/B7 , \picorv32_core/pcpi_rs2$25$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b25/or_B0_B1  (\picorv32_core/sel42_b25/or_B0_B1_o , \picorv32_core/sel42_b25/B0 , \picorv32_core/sel42_b25/B1 );
  or \picorv32_core/sel42_b25/or_B2_B3  (\picorv32_core/sel42_b25/or_B2_B3_o , \picorv32_core/sel42_b25/B2 , \picorv32_core/sel42_b25/B3 );
  or \picorv32_core/sel42_b25/or_B4_B5  (\picorv32_core/sel42_b25/or_B4_B5_o , \picorv32_core/sel42_b25/B4 , \picorv32_core/sel42_b25/B5 );
  or \picorv32_core/sel42_b25/or_B6_B7  (\picorv32_core/sel42_b25/or_B6_B7_o , \picorv32_core/sel42_b25/B6 , \picorv32_core/sel42_b25/B7 );
  or \picorv32_core/sel42_b25/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b25/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b25/or_B0_B1_o , \picorv32_core/sel42_b25/or_B2_B3_o );
  or \picorv32_core/sel42_b25/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b25/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b25/or_B4_B5_o , \picorv32_core/sel42_b25/or_B6_B7_o );
  or \picorv32_core/sel42_b25/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [25], \picorv32_core/sel42_b25/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b25/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b26/and_b0_0  (\picorv32_core/sel42_b26/B0 , \picorv32_core/pcpi_rs2$26$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b26/and_b0_1  (\picorv32_core/sel42_b26/B1 , \picorv32_core/pcpi_rs2$26$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b26/and_b0_2  (\picorv32_core/sel42_b26/B2 , \picorv32_core/pcpi_rs2$26$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b26/and_b0_3  (\picorv32_core/sel42_b26/B3 , \picorv32_core/pcpi_rs2$26$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b26/and_b0_4  (\picorv32_core/sel42_b26/B4 , \picorv32_core/cpuregs_rs2 [26], \picorv32_core/n665 );
  and \picorv32_core/sel42_b26/and_b0_5  (\picorv32_core/sel42_b26/B5 , \picorv32_core/n528 [26], \picorv32_core/n664 );
  and \picorv32_core/sel42_b26/and_b0_6  (\picorv32_core/sel42_b26/B6 , \picorv32_core/pcpi_rs2$26$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b26/and_b0_7  (\picorv32_core/sel42_b26/B7 , \picorv32_core/pcpi_rs2$26$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b26/or_B0_B1  (\picorv32_core/sel42_b26/or_B0_B1_o , \picorv32_core/sel42_b26/B0 , \picorv32_core/sel42_b26/B1 );
  or \picorv32_core/sel42_b26/or_B2_B3  (\picorv32_core/sel42_b26/or_B2_B3_o , \picorv32_core/sel42_b26/B2 , \picorv32_core/sel42_b26/B3 );
  or \picorv32_core/sel42_b26/or_B4_B5  (\picorv32_core/sel42_b26/or_B4_B5_o , \picorv32_core/sel42_b26/B4 , \picorv32_core/sel42_b26/B5 );
  or \picorv32_core/sel42_b26/or_B6_B7  (\picorv32_core/sel42_b26/or_B6_B7_o , \picorv32_core/sel42_b26/B6 , \picorv32_core/sel42_b26/B7 );
  or \picorv32_core/sel42_b26/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b26/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b26/or_B0_B1_o , \picorv32_core/sel42_b26/or_B2_B3_o );
  or \picorv32_core/sel42_b26/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b26/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b26/or_B4_B5_o , \picorv32_core/sel42_b26/or_B6_B7_o );
  or \picorv32_core/sel42_b26/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [26], \picorv32_core/sel42_b26/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b26/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b27/and_b0_0  (\picorv32_core/sel42_b27/B0 , \picorv32_core/pcpi_rs2$27$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b27/and_b0_1  (\picorv32_core/sel42_b27/B1 , \picorv32_core/pcpi_rs2$27$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b27/and_b0_2  (\picorv32_core/sel42_b27/B2 , \picorv32_core/pcpi_rs2$27$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b27/and_b0_3  (\picorv32_core/sel42_b27/B3 , \picorv32_core/pcpi_rs2$27$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b27/and_b0_4  (\picorv32_core/sel42_b27/B4 , \picorv32_core/cpuregs_rs2 [27], \picorv32_core/n665 );
  and \picorv32_core/sel42_b27/and_b0_5  (\picorv32_core/sel42_b27/B5 , \picorv32_core/n528 [27], \picorv32_core/n664 );
  and \picorv32_core/sel42_b27/and_b0_6  (\picorv32_core/sel42_b27/B6 , \picorv32_core/pcpi_rs2$27$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b27/and_b0_7  (\picorv32_core/sel42_b27/B7 , \picorv32_core/pcpi_rs2$27$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b27/or_B0_B1  (\picorv32_core/sel42_b27/or_B0_B1_o , \picorv32_core/sel42_b27/B0 , \picorv32_core/sel42_b27/B1 );
  or \picorv32_core/sel42_b27/or_B2_B3  (\picorv32_core/sel42_b27/or_B2_B3_o , \picorv32_core/sel42_b27/B2 , \picorv32_core/sel42_b27/B3 );
  or \picorv32_core/sel42_b27/or_B4_B5  (\picorv32_core/sel42_b27/or_B4_B5_o , \picorv32_core/sel42_b27/B4 , \picorv32_core/sel42_b27/B5 );
  or \picorv32_core/sel42_b27/or_B6_B7  (\picorv32_core/sel42_b27/or_B6_B7_o , \picorv32_core/sel42_b27/B6 , \picorv32_core/sel42_b27/B7 );
  or \picorv32_core/sel42_b27/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b27/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b27/or_B0_B1_o , \picorv32_core/sel42_b27/or_B2_B3_o );
  or \picorv32_core/sel42_b27/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b27/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b27/or_B4_B5_o , \picorv32_core/sel42_b27/or_B6_B7_o );
  or \picorv32_core/sel42_b27/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [27], \picorv32_core/sel42_b27/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b27/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b28/and_b0_0  (\picorv32_core/sel42_b28/B0 , \picorv32_core/pcpi_rs2$28$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b28/and_b0_1  (\picorv32_core/sel42_b28/B1 , \picorv32_core/pcpi_rs2$28$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b28/and_b0_2  (\picorv32_core/sel42_b28/B2 , \picorv32_core/pcpi_rs2$28$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b28/and_b0_3  (\picorv32_core/sel42_b28/B3 , \picorv32_core/pcpi_rs2$28$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b28/and_b0_4  (\picorv32_core/sel42_b28/B4 , \picorv32_core/cpuregs_rs2 [28], \picorv32_core/n665 );
  and \picorv32_core/sel42_b28/and_b0_5  (\picorv32_core/sel42_b28/B5 , \picorv32_core/n528 [28], \picorv32_core/n664 );
  and \picorv32_core/sel42_b28/and_b0_6  (\picorv32_core/sel42_b28/B6 , \picorv32_core/pcpi_rs2$28$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b28/and_b0_7  (\picorv32_core/sel42_b28/B7 , \picorv32_core/pcpi_rs2$28$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b28/or_B0_B1  (\picorv32_core/sel42_b28/or_B0_B1_o , \picorv32_core/sel42_b28/B0 , \picorv32_core/sel42_b28/B1 );
  or \picorv32_core/sel42_b28/or_B2_B3  (\picorv32_core/sel42_b28/or_B2_B3_o , \picorv32_core/sel42_b28/B2 , \picorv32_core/sel42_b28/B3 );
  or \picorv32_core/sel42_b28/or_B4_B5  (\picorv32_core/sel42_b28/or_B4_B5_o , \picorv32_core/sel42_b28/B4 , \picorv32_core/sel42_b28/B5 );
  or \picorv32_core/sel42_b28/or_B6_B7  (\picorv32_core/sel42_b28/or_B6_B7_o , \picorv32_core/sel42_b28/B6 , \picorv32_core/sel42_b28/B7 );
  or \picorv32_core/sel42_b28/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b28/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b28/or_B0_B1_o , \picorv32_core/sel42_b28/or_B2_B3_o );
  or \picorv32_core/sel42_b28/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b28/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b28/or_B4_B5_o , \picorv32_core/sel42_b28/or_B6_B7_o );
  or \picorv32_core/sel42_b28/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [28], \picorv32_core/sel42_b28/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b28/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b29/and_b0_0  (\picorv32_core/sel42_b29/B0 , \picorv32_core/pcpi_rs2$29$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b29/and_b0_1  (\picorv32_core/sel42_b29/B1 , \picorv32_core/pcpi_rs2$29$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b29/and_b0_2  (\picorv32_core/sel42_b29/B2 , \picorv32_core/pcpi_rs2$29$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b29/and_b0_3  (\picorv32_core/sel42_b29/B3 , \picorv32_core/pcpi_rs2$29$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b29/and_b0_4  (\picorv32_core/sel42_b29/B4 , \picorv32_core/cpuregs_rs2 [29], \picorv32_core/n665 );
  and \picorv32_core/sel42_b29/and_b0_5  (\picorv32_core/sel42_b29/B5 , \picorv32_core/n528 [29], \picorv32_core/n664 );
  and \picorv32_core/sel42_b29/and_b0_6  (\picorv32_core/sel42_b29/B6 , \picorv32_core/pcpi_rs2$29$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b29/and_b0_7  (\picorv32_core/sel42_b29/B7 , \picorv32_core/pcpi_rs2$29$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b29/or_B0_B1  (\picorv32_core/sel42_b29/or_B0_B1_o , \picorv32_core/sel42_b29/B0 , \picorv32_core/sel42_b29/B1 );
  or \picorv32_core/sel42_b29/or_B2_B3  (\picorv32_core/sel42_b29/or_B2_B3_o , \picorv32_core/sel42_b29/B2 , \picorv32_core/sel42_b29/B3 );
  or \picorv32_core/sel42_b29/or_B4_B5  (\picorv32_core/sel42_b29/or_B4_B5_o , \picorv32_core/sel42_b29/B4 , \picorv32_core/sel42_b29/B5 );
  or \picorv32_core/sel42_b29/or_B6_B7  (\picorv32_core/sel42_b29/or_B6_B7_o , \picorv32_core/sel42_b29/B6 , \picorv32_core/sel42_b29/B7 );
  or \picorv32_core/sel42_b29/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b29/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b29/or_B0_B1_o , \picorv32_core/sel42_b29/or_B2_B3_o );
  or \picorv32_core/sel42_b29/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b29/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b29/or_B4_B5_o , \picorv32_core/sel42_b29/or_B6_B7_o );
  or \picorv32_core/sel42_b29/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [29], \picorv32_core/sel42_b29/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b29/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b3/and_b0_0  (\picorv32_core/sel42_b3/B0 , mem_la_wdata[3], \picorv32_core/n669 );
  and \picorv32_core/sel42_b3/and_b0_1  (\picorv32_core/sel42_b3/B1 , mem_la_wdata[3], \picorv32_core/n668 );
  and \picorv32_core/sel42_b3/and_b0_2  (\picorv32_core/sel42_b3/B2 , mem_la_wdata[3], \picorv32_core/n667 );
  and \picorv32_core/sel42_b3/and_b0_3  (\picorv32_core/sel42_b3/B3 , mem_la_wdata[3], \picorv32_core/n666 );
  and \picorv32_core/sel42_b3/and_b0_4  (\picorv32_core/sel42_b3/B4 , \picorv32_core/cpuregs_rs2 [3], \picorv32_core/n665 );
  and \picorv32_core/sel42_b3/and_b0_5  (\picorv32_core/sel42_b3/B5 , \picorv32_core/n528 [3], \picorv32_core/n664 );
  and \picorv32_core/sel42_b3/and_b0_6  (\picorv32_core/sel42_b3/B6 , mem_la_wdata[3], \picorv32_core/n663 );
  and \picorv32_core/sel42_b3/and_b0_7  (\picorv32_core/sel42_b3/B7 , mem_la_wdata[3], \picorv32_core/n662 );
  or \picorv32_core/sel42_b3/or_B0_B1  (\picorv32_core/sel42_b3/or_B0_B1_o , \picorv32_core/sel42_b3/B0 , \picorv32_core/sel42_b3/B1 );
  or \picorv32_core/sel42_b3/or_B2_B3  (\picorv32_core/sel42_b3/or_B2_B3_o , \picorv32_core/sel42_b3/B2 , \picorv32_core/sel42_b3/B3 );
  or \picorv32_core/sel42_b3/or_B4_B5  (\picorv32_core/sel42_b3/or_B4_B5_o , \picorv32_core/sel42_b3/B4 , \picorv32_core/sel42_b3/B5 );
  or \picorv32_core/sel42_b3/or_B6_B7  (\picorv32_core/sel42_b3/or_B6_B7_o , \picorv32_core/sel42_b3/B6 , \picorv32_core/sel42_b3/B7 );
  or \picorv32_core/sel42_b3/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b3/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b3/or_B0_B1_o , \picorv32_core/sel42_b3/or_B2_B3_o );
  or \picorv32_core/sel42_b3/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b3/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b3/or_B4_B5_o , \picorv32_core/sel42_b3/or_B6_B7_o );
  or \picorv32_core/sel42_b3/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [3], \picorv32_core/sel42_b3/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b3/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b30/and_b0_0  (\picorv32_core/sel42_b30/B0 , \picorv32_core/pcpi_rs2$30$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b30/and_b0_1  (\picorv32_core/sel42_b30/B1 , \picorv32_core/pcpi_rs2$30$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b30/and_b0_2  (\picorv32_core/sel42_b30/B2 , \picorv32_core/pcpi_rs2$30$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b30/and_b0_3  (\picorv32_core/sel42_b30/B3 , \picorv32_core/pcpi_rs2$30$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b30/and_b0_4  (\picorv32_core/sel42_b30/B4 , \picorv32_core/cpuregs_rs2 [30], \picorv32_core/n665 );
  and \picorv32_core/sel42_b30/and_b0_5  (\picorv32_core/sel42_b30/B5 , \picorv32_core/n528 [30], \picorv32_core/n664 );
  and \picorv32_core/sel42_b30/and_b0_6  (\picorv32_core/sel42_b30/B6 , \picorv32_core/pcpi_rs2$30$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b30/and_b0_7  (\picorv32_core/sel42_b30/B7 , \picorv32_core/pcpi_rs2$30$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b30/or_B0_B1  (\picorv32_core/sel42_b30/or_B0_B1_o , \picorv32_core/sel42_b30/B0 , \picorv32_core/sel42_b30/B1 );
  or \picorv32_core/sel42_b30/or_B2_B3  (\picorv32_core/sel42_b30/or_B2_B3_o , \picorv32_core/sel42_b30/B2 , \picorv32_core/sel42_b30/B3 );
  or \picorv32_core/sel42_b30/or_B4_B5  (\picorv32_core/sel42_b30/or_B4_B5_o , \picorv32_core/sel42_b30/B4 , \picorv32_core/sel42_b30/B5 );
  or \picorv32_core/sel42_b30/or_B6_B7  (\picorv32_core/sel42_b30/or_B6_B7_o , \picorv32_core/sel42_b30/B6 , \picorv32_core/sel42_b30/B7 );
  or \picorv32_core/sel42_b30/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b30/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b30/or_B0_B1_o , \picorv32_core/sel42_b30/or_B2_B3_o );
  or \picorv32_core/sel42_b30/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b30/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b30/or_B4_B5_o , \picorv32_core/sel42_b30/or_B6_B7_o );
  or \picorv32_core/sel42_b30/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [30], \picorv32_core/sel42_b30/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b30/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b31/and_b0_0  (\picorv32_core/sel42_b31/B0 , \picorv32_core/pcpi_rs2$31$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b31/and_b0_1  (\picorv32_core/sel42_b31/B1 , \picorv32_core/pcpi_rs2$31$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b31/and_b0_2  (\picorv32_core/sel42_b31/B2 , \picorv32_core/pcpi_rs2$31$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b31/and_b0_3  (\picorv32_core/sel42_b31/B3 , \picorv32_core/pcpi_rs2$31$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b31/and_b0_4  (\picorv32_core/sel42_b31/B4 , \picorv32_core/cpuregs_rs2 [31], \picorv32_core/n665 );
  and \picorv32_core/sel42_b31/and_b0_5  (\picorv32_core/sel42_b31/B5 , \picorv32_core/n528 [31], \picorv32_core/n664 );
  and \picorv32_core/sel42_b31/and_b0_6  (\picorv32_core/sel42_b31/B6 , \picorv32_core/pcpi_rs2$31$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b31/and_b0_7  (\picorv32_core/sel42_b31/B7 , \picorv32_core/pcpi_rs2$31$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b31/or_B0_B1  (\picorv32_core/sel42_b31/or_B0_B1_o , \picorv32_core/sel42_b31/B0 , \picorv32_core/sel42_b31/B1 );
  or \picorv32_core/sel42_b31/or_B2_B3  (\picorv32_core/sel42_b31/or_B2_B3_o , \picorv32_core/sel42_b31/B2 , \picorv32_core/sel42_b31/B3 );
  or \picorv32_core/sel42_b31/or_B4_B5  (\picorv32_core/sel42_b31/or_B4_B5_o , \picorv32_core/sel42_b31/B4 , \picorv32_core/sel42_b31/B5 );
  or \picorv32_core/sel42_b31/or_B6_B7  (\picorv32_core/sel42_b31/or_B6_B7_o , \picorv32_core/sel42_b31/B6 , \picorv32_core/sel42_b31/B7 );
  or \picorv32_core/sel42_b31/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b31/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b31/or_B0_B1_o , \picorv32_core/sel42_b31/or_B2_B3_o );
  or \picorv32_core/sel42_b31/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b31/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b31/or_B4_B5_o , \picorv32_core/sel42_b31/or_B6_B7_o );
  or \picorv32_core/sel42_b31/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [31], \picorv32_core/sel42_b31/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b31/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b4/and_b0_0  (\picorv32_core/sel42_b4/B0 , mem_la_wdata[4], \picorv32_core/n669 );
  and \picorv32_core/sel42_b4/and_b0_1  (\picorv32_core/sel42_b4/B1 , mem_la_wdata[4], \picorv32_core/n668 );
  and \picorv32_core/sel42_b4/and_b0_2  (\picorv32_core/sel42_b4/B2 , mem_la_wdata[4], \picorv32_core/n667 );
  and \picorv32_core/sel42_b4/and_b0_3  (\picorv32_core/sel42_b4/B3 , mem_la_wdata[4], \picorv32_core/n666 );
  and \picorv32_core/sel42_b4/and_b0_4  (\picorv32_core/sel42_b4/B4 , \picorv32_core/cpuregs_rs2 [4], \picorv32_core/n665 );
  and \picorv32_core/sel42_b4/and_b0_5  (\picorv32_core/sel42_b4/B5 , \picorv32_core/n528 [4], \picorv32_core/n664 );
  and \picorv32_core/sel42_b4/and_b0_6  (\picorv32_core/sel42_b4/B6 , mem_la_wdata[4], \picorv32_core/n663 );
  and \picorv32_core/sel42_b4/and_b0_7  (\picorv32_core/sel42_b4/B7 , mem_la_wdata[4], \picorv32_core/n662 );
  or \picorv32_core/sel42_b4/or_B0_B1  (\picorv32_core/sel42_b4/or_B0_B1_o , \picorv32_core/sel42_b4/B0 , \picorv32_core/sel42_b4/B1 );
  or \picorv32_core/sel42_b4/or_B2_B3  (\picorv32_core/sel42_b4/or_B2_B3_o , \picorv32_core/sel42_b4/B2 , \picorv32_core/sel42_b4/B3 );
  or \picorv32_core/sel42_b4/or_B4_B5  (\picorv32_core/sel42_b4/or_B4_B5_o , \picorv32_core/sel42_b4/B4 , \picorv32_core/sel42_b4/B5 );
  or \picorv32_core/sel42_b4/or_B6_B7  (\picorv32_core/sel42_b4/or_B6_B7_o , \picorv32_core/sel42_b4/B6 , \picorv32_core/sel42_b4/B7 );
  or \picorv32_core/sel42_b4/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b4/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b4/or_B0_B1_o , \picorv32_core/sel42_b4/or_B2_B3_o );
  or \picorv32_core/sel42_b4/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b4/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b4/or_B4_B5_o , \picorv32_core/sel42_b4/or_B6_B7_o );
  or \picorv32_core/sel42_b4/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [4], \picorv32_core/sel42_b4/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b4/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b5/and_b0_0  (\picorv32_core/sel42_b5/B0 , mem_la_wdata[5], \picorv32_core/n669 );
  and \picorv32_core/sel42_b5/and_b0_1  (\picorv32_core/sel42_b5/B1 , mem_la_wdata[5], \picorv32_core/n668 );
  and \picorv32_core/sel42_b5/and_b0_2  (\picorv32_core/sel42_b5/B2 , mem_la_wdata[5], \picorv32_core/n667 );
  and \picorv32_core/sel42_b5/and_b0_3  (\picorv32_core/sel42_b5/B3 , mem_la_wdata[5], \picorv32_core/n666 );
  and \picorv32_core/sel42_b5/and_b0_4  (\picorv32_core/sel42_b5/B4 , \picorv32_core/cpuregs_rs2 [5], \picorv32_core/n665 );
  and \picorv32_core/sel42_b5/and_b0_5  (\picorv32_core/sel42_b5/B5 , \picorv32_core/n528 [5], \picorv32_core/n664 );
  and \picorv32_core/sel42_b5/and_b0_6  (\picorv32_core/sel42_b5/B6 , mem_la_wdata[5], \picorv32_core/n663 );
  and \picorv32_core/sel42_b5/and_b0_7  (\picorv32_core/sel42_b5/B7 , mem_la_wdata[5], \picorv32_core/n662 );
  or \picorv32_core/sel42_b5/or_B0_B1  (\picorv32_core/sel42_b5/or_B0_B1_o , \picorv32_core/sel42_b5/B0 , \picorv32_core/sel42_b5/B1 );
  or \picorv32_core/sel42_b5/or_B2_B3  (\picorv32_core/sel42_b5/or_B2_B3_o , \picorv32_core/sel42_b5/B2 , \picorv32_core/sel42_b5/B3 );
  or \picorv32_core/sel42_b5/or_B4_B5  (\picorv32_core/sel42_b5/or_B4_B5_o , \picorv32_core/sel42_b5/B4 , \picorv32_core/sel42_b5/B5 );
  or \picorv32_core/sel42_b5/or_B6_B7  (\picorv32_core/sel42_b5/or_B6_B7_o , \picorv32_core/sel42_b5/B6 , \picorv32_core/sel42_b5/B7 );
  or \picorv32_core/sel42_b5/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b5/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b5/or_B0_B1_o , \picorv32_core/sel42_b5/or_B2_B3_o );
  or \picorv32_core/sel42_b5/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b5/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b5/or_B4_B5_o , \picorv32_core/sel42_b5/or_B6_B7_o );
  or \picorv32_core/sel42_b5/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [5], \picorv32_core/sel42_b5/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b5/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b6/and_b0_0  (\picorv32_core/sel42_b6/B0 , mem_la_wdata[6], \picorv32_core/n669 );
  and \picorv32_core/sel42_b6/and_b0_1  (\picorv32_core/sel42_b6/B1 , mem_la_wdata[6], \picorv32_core/n668 );
  and \picorv32_core/sel42_b6/and_b0_2  (\picorv32_core/sel42_b6/B2 , mem_la_wdata[6], \picorv32_core/n667 );
  and \picorv32_core/sel42_b6/and_b0_3  (\picorv32_core/sel42_b6/B3 , mem_la_wdata[6], \picorv32_core/n666 );
  and \picorv32_core/sel42_b6/and_b0_4  (\picorv32_core/sel42_b6/B4 , \picorv32_core/cpuregs_rs2 [6], \picorv32_core/n665 );
  and \picorv32_core/sel42_b6/and_b0_5  (\picorv32_core/sel42_b6/B5 , \picorv32_core/n528 [6], \picorv32_core/n664 );
  and \picorv32_core/sel42_b6/and_b0_6  (\picorv32_core/sel42_b6/B6 , mem_la_wdata[6], \picorv32_core/n663 );
  and \picorv32_core/sel42_b6/and_b0_7  (\picorv32_core/sel42_b6/B7 , mem_la_wdata[6], \picorv32_core/n662 );
  or \picorv32_core/sel42_b6/or_B0_B1  (\picorv32_core/sel42_b6/or_B0_B1_o , \picorv32_core/sel42_b6/B0 , \picorv32_core/sel42_b6/B1 );
  or \picorv32_core/sel42_b6/or_B2_B3  (\picorv32_core/sel42_b6/or_B2_B3_o , \picorv32_core/sel42_b6/B2 , \picorv32_core/sel42_b6/B3 );
  or \picorv32_core/sel42_b6/or_B4_B5  (\picorv32_core/sel42_b6/or_B4_B5_o , \picorv32_core/sel42_b6/B4 , \picorv32_core/sel42_b6/B5 );
  or \picorv32_core/sel42_b6/or_B6_B7  (\picorv32_core/sel42_b6/or_B6_B7_o , \picorv32_core/sel42_b6/B6 , \picorv32_core/sel42_b6/B7 );
  or \picorv32_core/sel42_b6/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b6/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b6/or_B0_B1_o , \picorv32_core/sel42_b6/or_B2_B3_o );
  or \picorv32_core/sel42_b6/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b6/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b6/or_B4_B5_o , \picorv32_core/sel42_b6/or_B6_B7_o );
  or \picorv32_core/sel42_b6/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [6], \picorv32_core/sel42_b6/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b6/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b7/and_b0_0  (\picorv32_core/sel42_b7/B0 , mem_la_wdata[7], \picorv32_core/n669 );
  and \picorv32_core/sel42_b7/and_b0_1  (\picorv32_core/sel42_b7/B1 , mem_la_wdata[7], \picorv32_core/n668 );
  and \picorv32_core/sel42_b7/and_b0_2  (\picorv32_core/sel42_b7/B2 , mem_la_wdata[7], \picorv32_core/n667 );
  and \picorv32_core/sel42_b7/and_b0_3  (\picorv32_core/sel42_b7/B3 , mem_la_wdata[7], \picorv32_core/n666 );
  and \picorv32_core/sel42_b7/and_b0_4  (\picorv32_core/sel42_b7/B4 , \picorv32_core/cpuregs_rs2 [7], \picorv32_core/n665 );
  and \picorv32_core/sel42_b7/and_b0_5  (\picorv32_core/sel42_b7/B5 , \picorv32_core/n528 [7], \picorv32_core/n664 );
  and \picorv32_core/sel42_b7/and_b0_6  (\picorv32_core/sel42_b7/B6 , mem_la_wdata[7], \picorv32_core/n663 );
  and \picorv32_core/sel42_b7/and_b0_7  (\picorv32_core/sel42_b7/B7 , mem_la_wdata[7], \picorv32_core/n662 );
  or \picorv32_core/sel42_b7/or_B0_B1  (\picorv32_core/sel42_b7/or_B0_B1_o , \picorv32_core/sel42_b7/B0 , \picorv32_core/sel42_b7/B1 );
  or \picorv32_core/sel42_b7/or_B2_B3  (\picorv32_core/sel42_b7/or_B2_B3_o , \picorv32_core/sel42_b7/B2 , \picorv32_core/sel42_b7/B3 );
  or \picorv32_core/sel42_b7/or_B4_B5  (\picorv32_core/sel42_b7/or_B4_B5_o , \picorv32_core/sel42_b7/B4 , \picorv32_core/sel42_b7/B5 );
  or \picorv32_core/sel42_b7/or_B6_B7  (\picorv32_core/sel42_b7/or_B6_B7_o , \picorv32_core/sel42_b7/B6 , \picorv32_core/sel42_b7/B7 );
  or \picorv32_core/sel42_b7/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b7/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b7/or_B0_B1_o , \picorv32_core/sel42_b7/or_B2_B3_o );
  or \picorv32_core/sel42_b7/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b7/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b7/or_B4_B5_o , \picorv32_core/sel42_b7/or_B6_B7_o );
  or \picorv32_core/sel42_b7/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [7], \picorv32_core/sel42_b7/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b7/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b8/and_b0_0  (\picorv32_core/sel42_b8/B0 , \picorv32_core/pcpi_rs2$8$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b8/and_b0_1  (\picorv32_core/sel42_b8/B1 , \picorv32_core/pcpi_rs2$8$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b8/and_b0_2  (\picorv32_core/sel42_b8/B2 , \picorv32_core/pcpi_rs2$8$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b8/and_b0_3  (\picorv32_core/sel42_b8/B3 , \picorv32_core/pcpi_rs2$8$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b8/and_b0_4  (\picorv32_core/sel42_b8/B4 , \picorv32_core/cpuregs_rs2 [8], \picorv32_core/n665 );
  and \picorv32_core/sel42_b8/and_b0_5  (\picorv32_core/sel42_b8/B5 , \picorv32_core/n528 [8], \picorv32_core/n664 );
  and \picorv32_core/sel42_b8/and_b0_6  (\picorv32_core/sel42_b8/B6 , \picorv32_core/pcpi_rs2$8$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b8/and_b0_7  (\picorv32_core/sel42_b8/B7 , \picorv32_core/pcpi_rs2$8$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b8/or_B0_B1  (\picorv32_core/sel42_b8/or_B0_B1_o , \picorv32_core/sel42_b8/B0 , \picorv32_core/sel42_b8/B1 );
  or \picorv32_core/sel42_b8/or_B2_B3  (\picorv32_core/sel42_b8/or_B2_B3_o , \picorv32_core/sel42_b8/B2 , \picorv32_core/sel42_b8/B3 );
  or \picorv32_core/sel42_b8/or_B4_B5  (\picorv32_core/sel42_b8/or_B4_B5_o , \picorv32_core/sel42_b8/B4 , \picorv32_core/sel42_b8/B5 );
  or \picorv32_core/sel42_b8/or_B6_B7  (\picorv32_core/sel42_b8/or_B6_B7_o , \picorv32_core/sel42_b8/B6 , \picorv32_core/sel42_b8/B7 );
  or \picorv32_core/sel42_b8/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b8/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b8/or_B0_B1_o , \picorv32_core/sel42_b8/or_B2_B3_o );
  or \picorv32_core/sel42_b8/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b8/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b8/or_B4_B5_o , \picorv32_core/sel42_b8/or_B6_B7_o );
  or \picorv32_core/sel42_b8/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [8], \picorv32_core/sel42_b8/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b8/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel42_b9/and_b0_0  (\picorv32_core/sel42_b9/B0 , \picorv32_core/pcpi_rs2$9$ , \picorv32_core/n669 );
  and \picorv32_core/sel42_b9/and_b0_1  (\picorv32_core/sel42_b9/B1 , \picorv32_core/pcpi_rs2$9$ , \picorv32_core/n668 );
  and \picorv32_core/sel42_b9/and_b0_2  (\picorv32_core/sel42_b9/B2 , \picorv32_core/pcpi_rs2$9$ , \picorv32_core/n667 );
  and \picorv32_core/sel42_b9/and_b0_3  (\picorv32_core/sel42_b9/B3 , \picorv32_core/pcpi_rs2$9$ , \picorv32_core/n666 );
  and \picorv32_core/sel42_b9/and_b0_4  (\picorv32_core/sel42_b9/B4 , \picorv32_core/cpuregs_rs2 [9], \picorv32_core/n665 );
  and \picorv32_core/sel42_b9/and_b0_5  (\picorv32_core/sel42_b9/B5 , \picorv32_core/n528 [9], \picorv32_core/n664 );
  and \picorv32_core/sel42_b9/and_b0_6  (\picorv32_core/sel42_b9/B6 , \picorv32_core/pcpi_rs2$9$ , \picorv32_core/n663 );
  and \picorv32_core/sel42_b9/and_b0_7  (\picorv32_core/sel42_b9/B7 , \picorv32_core/pcpi_rs2$9$ , \picorv32_core/n662 );
  or \picorv32_core/sel42_b9/or_B0_B1  (\picorv32_core/sel42_b9/or_B0_B1_o , \picorv32_core/sel42_b9/B0 , \picorv32_core/sel42_b9/B1 );
  or \picorv32_core/sel42_b9/or_B2_B3  (\picorv32_core/sel42_b9/or_B2_B3_o , \picorv32_core/sel42_b9/B2 , \picorv32_core/sel42_b9/B3 );
  or \picorv32_core/sel42_b9/or_B4_B5  (\picorv32_core/sel42_b9/or_B4_B5_o , \picorv32_core/sel42_b9/B4 , \picorv32_core/sel42_b9/B5 );
  or \picorv32_core/sel42_b9/or_B6_B7  (\picorv32_core/sel42_b9/or_B6_B7_o , \picorv32_core/sel42_b9/B6 , \picorv32_core/sel42_b9/B7 );
  or \picorv32_core/sel42_b9/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel42_b9/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b9/or_B0_B1_o , \picorv32_core/sel42_b9/or_B2_B3_o );
  or \picorv32_core/sel42_b9/or_or_B4_B5_o_or_B6_  (\picorv32_core/sel42_b9/or_or_B4_B5_o_or_B6__o , \picorv32_core/sel42_b9/or_B4_B5_o , \picorv32_core/sel42_b9/or_B6_B7_o );
  or \picorv32_core/sel42_b9/or_or_or_B0_B1_o_or_  (\picorv32_core/n694 [9], \picorv32_core/sel42_b9/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel42_b9/or_or_B4_B5_o_or_B6__o );
  and \picorv32_core/sel43_b0/and_b0_0  (\picorv32_core/sel43_b0/B0 , \picorv32_core/n658 [0], \picorv32_core/n669 );
  and \picorv32_core/sel43_b0/and_b0_2  (\picorv32_core/sel43_b0/B2 , \picorv32_core/n567 [0], \picorv32_core/n667 );
  and \picorv32_core/sel43_b0/and_b0_3  (\picorv32_core/sel43_b0/B3 , \picorv32_core/n543 [0], \picorv32_core/n666 );
  and \picorv32_core/sel43_b0/and_b0_5  (\picorv32_core/sel43_b0/B5 , \picorv32_core/n525 [0], \picorv32_core/n664 );
  or \picorv32_core/sel43_b0/or_B2_B3  (\picorv32_core/sel43_b0/or_B2_B3_o , \picorv32_core/sel43_b0/B2 , \picorv32_core/sel43_b0/B3 );
  or \picorv32_core/sel43_b0/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b0/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b0/B0 , \picorv32_core/sel43_b0/or_B2_B3_o );
  or \picorv32_core/sel43_b0/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [0], \picorv32_core/sel43_b0/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b0/B5 );
  and \picorv32_core/sel43_b1/and_b0_0  (\picorv32_core/sel43_b1/B0 , \picorv32_core/n658 [1], \picorv32_core/n669 );
  and \picorv32_core/sel43_b1/and_b0_2  (\picorv32_core/sel43_b1/B2 , \picorv32_core/n567 [1], \picorv32_core/n667 );
  and \picorv32_core/sel43_b1/and_b0_3  (\picorv32_core/sel43_b1/B3 , \picorv32_core/n543 [1], \picorv32_core/n666 );
  and \picorv32_core/sel43_b1/and_b0_5  (\picorv32_core/sel43_b1/B5 , \picorv32_core/n525 [1], \picorv32_core/n664 );
  or \picorv32_core/sel43_b1/or_B2_B3  (\picorv32_core/sel43_b1/or_B2_B3_o , \picorv32_core/sel43_b1/B2 , \picorv32_core/sel43_b1/B3 );
  or \picorv32_core/sel43_b1/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b1/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b1/B0 , \picorv32_core/sel43_b1/or_B2_B3_o );
  or \picorv32_core/sel43_b1/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [1], \picorv32_core/sel43_b1/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b1/B5 );
  and \picorv32_core/sel43_b10/and_b0_0  (\picorv32_core/sel43_b10/B0 , \picorv32_core/n658 [10], \picorv32_core/n669 );
  and \picorv32_core/sel43_b10/and_b0_2  (\picorv32_core/sel43_b10/B2 , \picorv32_core/n567 [10], \picorv32_core/n667 );
  and \picorv32_core/sel43_b10/and_b0_3  (\picorv32_core/sel43_b10/B3 , \picorv32_core/n543 [10], \picorv32_core/n666 );
  and \picorv32_core/sel43_b10/and_b0_5  (\picorv32_core/sel43_b10/B5 , \picorv32_core/n525 [10], \picorv32_core/n664 );
  or \picorv32_core/sel43_b10/or_B2_B3  (\picorv32_core/sel43_b10/or_B2_B3_o , \picorv32_core/sel43_b10/B2 , \picorv32_core/sel43_b10/B3 );
  or \picorv32_core/sel43_b10/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b10/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b10/B0 , \picorv32_core/sel43_b10/or_B2_B3_o );
  or \picorv32_core/sel43_b10/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [10], \picorv32_core/sel43_b10/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b10/B5 );
  and \picorv32_core/sel43_b11/and_b0_0  (\picorv32_core/sel43_b11/B0 , \picorv32_core/n658 [11], \picorv32_core/n669 );
  and \picorv32_core/sel43_b11/and_b0_2  (\picorv32_core/sel43_b11/B2 , \picorv32_core/n567 [11], \picorv32_core/n667 );
  and \picorv32_core/sel43_b11/and_b0_3  (\picorv32_core/sel43_b11/B3 , \picorv32_core/n543 [11], \picorv32_core/n666 );
  and \picorv32_core/sel43_b11/and_b0_5  (\picorv32_core/sel43_b11/B5 , \picorv32_core/n525 [11], \picorv32_core/n664 );
  or \picorv32_core/sel43_b11/or_B2_B3  (\picorv32_core/sel43_b11/or_B2_B3_o , \picorv32_core/sel43_b11/B2 , \picorv32_core/sel43_b11/B3 );
  or \picorv32_core/sel43_b11/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b11/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b11/B0 , \picorv32_core/sel43_b11/or_B2_B3_o );
  or \picorv32_core/sel43_b11/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [11], \picorv32_core/sel43_b11/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b11/B5 );
  and \picorv32_core/sel43_b12/and_b0_0  (\picorv32_core/sel43_b12/B0 , \picorv32_core/n658 [12], \picorv32_core/n669 );
  and \picorv32_core/sel43_b12/and_b0_2  (\picorv32_core/sel43_b12/B2 , \picorv32_core/n567 [12], \picorv32_core/n667 );
  and \picorv32_core/sel43_b12/and_b0_3  (\picorv32_core/sel43_b12/B3 , \picorv32_core/n543 [12], \picorv32_core/n666 );
  and \picorv32_core/sel43_b12/and_b0_5  (\picorv32_core/sel43_b12/B5 , \picorv32_core/n525 [12], \picorv32_core/n664 );
  or \picorv32_core/sel43_b12/or_B2_B3  (\picorv32_core/sel43_b12/or_B2_B3_o , \picorv32_core/sel43_b12/B2 , \picorv32_core/sel43_b12/B3 );
  or \picorv32_core/sel43_b12/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b12/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b12/B0 , \picorv32_core/sel43_b12/or_B2_B3_o );
  or \picorv32_core/sel43_b12/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [12], \picorv32_core/sel43_b12/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b12/B5 );
  and \picorv32_core/sel43_b13/and_b0_0  (\picorv32_core/sel43_b13/B0 , \picorv32_core/n658 [13], \picorv32_core/n669 );
  and \picorv32_core/sel43_b13/and_b0_2  (\picorv32_core/sel43_b13/B2 , \picorv32_core/n567 [13], \picorv32_core/n667 );
  and \picorv32_core/sel43_b13/and_b0_3  (\picorv32_core/sel43_b13/B3 , \picorv32_core/n543 [13], \picorv32_core/n666 );
  and \picorv32_core/sel43_b13/and_b0_5  (\picorv32_core/sel43_b13/B5 , \picorv32_core/n525 [13], \picorv32_core/n664 );
  or \picorv32_core/sel43_b13/or_B2_B3  (\picorv32_core/sel43_b13/or_B2_B3_o , \picorv32_core/sel43_b13/B2 , \picorv32_core/sel43_b13/B3 );
  or \picorv32_core/sel43_b13/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b13/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b13/B0 , \picorv32_core/sel43_b13/or_B2_B3_o );
  or \picorv32_core/sel43_b13/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [13], \picorv32_core/sel43_b13/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b13/B5 );
  and \picorv32_core/sel43_b14/and_b0_0  (\picorv32_core/sel43_b14/B0 , \picorv32_core/n658 [14], \picorv32_core/n669 );
  and \picorv32_core/sel43_b14/and_b0_2  (\picorv32_core/sel43_b14/B2 , \picorv32_core/n567 [14], \picorv32_core/n667 );
  and \picorv32_core/sel43_b14/and_b0_3  (\picorv32_core/sel43_b14/B3 , \picorv32_core/n543 [14], \picorv32_core/n666 );
  and \picorv32_core/sel43_b14/and_b0_5  (\picorv32_core/sel43_b14/B5 , \picorv32_core/n525 [14], \picorv32_core/n664 );
  or \picorv32_core/sel43_b14/or_B2_B3  (\picorv32_core/sel43_b14/or_B2_B3_o , \picorv32_core/sel43_b14/B2 , \picorv32_core/sel43_b14/B3 );
  or \picorv32_core/sel43_b14/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b14/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b14/B0 , \picorv32_core/sel43_b14/or_B2_B3_o );
  or \picorv32_core/sel43_b14/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [14], \picorv32_core/sel43_b14/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b14/B5 );
  and \picorv32_core/sel43_b15/and_b0_0  (\picorv32_core/sel43_b15/B0 , \picorv32_core/n658 [15], \picorv32_core/n669 );
  and \picorv32_core/sel43_b15/and_b0_2  (\picorv32_core/sel43_b15/B2 , \picorv32_core/n567 [15], \picorv32_core/n667 );
  and \picorv32_core/sel43_b15/and_b0_3  (\picorv32_core/sel43_b15/B3 , \picorv32_core/n543 [15], \picorv32_core/n666 );
  and \picorv32_core/sel43_b15/and_b0_5  (\picorv32_core/sel43_b15/B5 , \picorv32_core/n525 [15], \picorv32_core/n664 );
  or \picorv32_core/sel43_b15/or_B2_B3  (\picorv32_core/sel43_b15/or_B2_B3_o , \picorv32_core/sel43_b15/B2 , \picorv32_core/sel43_b15/B3 );
  or \picorv32_core/sel43_b15/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b15/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b15/B0 , \picorv32_core/sel43_b15/or_B2_B3_o );
  or \picorv32_core/sel43_b15/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [15], \picorv32_core/sel43_b15/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b15/B5 );
  and \picorv32_core/sel43_b16/and_b0_0  (\picorv32_core/sel43_b16/B0 , \picorv32_core/n658 [16], \picorv32_core/n669 );
  and \picorv32_core/sel43_b16/and_b0_2  (\picorv32_core/sel43_b16/B2 , \picorv32_core/n567 [16], \picorv32_core/n667 );
  and \picorv32_core/sel43_b16/and_b0_3  (\picorv32_core/sel43_b16/B3 , \picorv32_core/n543 [16], \picorv32_core/n666 );
  and \picorv32_core/sel43_b16/and_b0_5  (\picorv32_core/sel43_b16/B5 , \picorv32_core/n525 [16], \picorv32_core/n664 );
  or \picorv32_core/sel43_b16/or_B2_B3  (\picorv32_core/sel43_b16/or_B2_B3_o , \picorv32_core/sel43_b16/B2 , \picorv32_core/sel43_b16/B3 );
  or \picorv32_core/sel43_b16/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b16/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b16/B0 , \picorv32_core/sel43_b16/or_B2_B3_o );
  or \picorv32_core/sel43_b16/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [16], \picorv32_core/sel43_b16/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b16/B5 );
  and \picorv32_core/sel43_b17/and_b0_0  (\picorv32_core/sel43_b17/B0 , \picorv32_core/n658 [17], \picorv32_core/n669 );
  and \picorv32_core/sel43_b17/and_b0_2  (\picorv32_core/sel43_b17/B2 , \picorv32_core/n567 [17], \picorv32_core/n667 );
  and \picorv32_core/sel43_b17/and_b0_3  (\picorv32_core/sel43_b17/B3 , \picorv32_core/n543 [17], \picorv32_core/n666 );
  and \picorv32_core/sel43_b17/and_b0_5  (\picorv32_core/sel43_b17/B5 , \picorv32_core/n525 [17], \picorv32_core/n664 );
  or \picorv32_core/sel43_b17/or_B2_B3  (\picorv32_core/sel43_b17/or_B2_B3_o , \picorv32_core/sel43_b17/B2 , \picorv32_core/sel43_b17/B3 );
  or \picorv32_core/sel43_b17/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b17/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b17/B0 , \picorv32_core/sel43_b17/or_B2_B3_o );
  or \picorv32_core/sel43_b17/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [17], \picorv32_core/sel43_b17/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b17/B5 );
  and \picorv32_core/sel43_b18/and_b0_0  (\picorv32_core/sel43_b18/B0 , \picorv32_core/n658 [18], \picorv32_core/n669 );
  and \picorv32_core/sel43_b18/and_b0_2  (\picorv32_core/sel43_b18/B2 , \picorv32_core/n567 [18], \picorv32_core/n667 );
  and \picorv32_core/sel43_b18/and_b0_3  (\picorv32_core/sel43_b18/B3 , \picorv32_core/n543 [18], \picorv32_core/n666 );
  and \picorv32_core/sel43_b18/and_b0_5  (\picorv32_core/sel43_b18/B5 , \picorv32_core/n525 [18], \picorv32_core/n664 );
  or \picorv32_core/sel43_b18/or_B2_B3  (\picorv32_core/sel43_b18/or_B2_B3_o , \picorv32_core/sel43_b18/B2 , \picorv32_core/sel43_b18/B3 );
  or \picorv32_core/sel43_b18/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b18/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b18/B0 , \picorv32_core/sel43_b18/or_B2_B3_o );
  or \picorv32_core/sel43_b18/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [18], \picorv32_core/sel43_b18/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b18/B5 );
  and \picorv32_core/sel43_b19/and_b0_0  (\picorv32_core/sel43_b19/B0 , \picorv32_core/n658 [19], \picorv32_core/n669 );
  and \picorv32_core/sel43_b19/and_b0_2  (\picorv32_core/sel43_b19/B2 , \picorv32_core/n567 [19], \picorv32_core/n667 );
  and \picorv32_core/sel43_b19/and_b0_3  (\picorv32_core/sel43_b19/B3 , \picorv32_core/n543 [19], \picorv32_core/n666 );
  and \picorv32_core/sel43_b19/and_b0_5  (\picorv32_core/sel43_b19/B5 , \picorv32_core/n525 [19], \picorv32_core/n664 );
  or \picorv32_core/sel43_b19/or_B2_B3  (\picorv32_core/sel43_b19/or_B2_B3_o , \picorv32_core/sel43_b19/B2 , \picorv32_core/sel43_b19/B3 );
  or \picorv32_core/sel43_b19/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b19/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b19/B0 , \picorv32_core/sel43_b19/or_B2_B3_o );
  or \picorv32_core/sel43_b19/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [19], \picorv32_core/sel43_b19/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b19/B5 );
  and \picorv32_core/sel43_b2/and_b0_0  (\picorv32_core/sel43_b2/B0 , \picorv32_core/n658 [2], \picorv32_core/n669 );
  and \picorv32_core/sel43_b2/and_b0_2  (\picorv32_core/sel43_b2/B2 , \picorv32_core/n567 [2], \picorv32_core/n667 );
  and \picorv32_core/sel43_b2/and_b0_3  (\picorv32_core/sel43_b2/B3 , \picorv32_core/n543 [2], \picorv32_core/n666 );
  and \picorv32_core/sel43_b2/and_b0_5  (\picorv32_core/sel43_b2/B5 , \picorv32_core/n525 [2], \picorv32_core/n664 );
  or \picorv32_core/sel43_b2/or_B2_B3  (\picorv32_core/sel43_b2/or_B2_B3_o , \picorv32_core/sel43_b2/B2 , \picorv32_core/sel43_b2/B3 );
  or \picorv32_core/sel43_b2/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b2/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b2/B0 , \picorv32_core/sel43_b2/or_B2_B3_o );
  or \picorv32_core/sel43_b2/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [2], \picorv32_core/sel43_b2/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b2/B5 );
  and \picorv32_core/sel43_b20/and_b0_0  (\picorv32_core/sel43_b20/B0 , \picorv32_core/n658 [20], \picorv32_core/n669 );
  and \picorv32_core/sel43_b20/and_b0_2  (\picorv32_core/sel43_b20/B2 , \picorv32_core/n567 [20], \picorv32_core/n667 );
  and \picorv32_core/sel43_b20/and_b0_3  (\picorv32_core/sel43_b20/B3 , \picorv32_core/n543 [20], \picorv32_core/n666 );
  and \picorv32_core/sel43_b20/and_b0_5  (\picorv32_core/sel43_b20/B5 , \picorv32_core/n525 [20], \picorv32_core/n664 );
  or \picorv32_core/sel43_b20/or_B2_B3  (\picorv32_core/sel43_b20/or_B2_B3_o , \picorv32_core/sel43_b20/B2 , \picorv32_core/sel43_b20/B3 );
  or \picorv32_core/sel43_b20/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b20/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b20/B0 , \picorv32_core/sel43_b20/or_B2_B3_o );
  or \picorv32_core/sel43_b20/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [20], \picorv32_core/sel43_b20/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b20/B5 );
  and \picorv32_core/sel43_b21/and_b0_0  (\picorv32_core/sel43_b21/B0 , \picorv32_core/n658 [21], \picorv32_core/n669 );
  and \picorv32_core/sel43_b21/and_b0_2  (\picorv32_core/sel43_b21/B2 , \picorv32_core/n567 [21], \picorv32_core/n667 );
  and \picorv32_core/sel43_b21/and_b0_3  (\picorv32_core/sel43_b21/B3 , \picorv32_core/n543 [21], \picorv32_core/n666 );
  and \picorv32_core/sel43_b21/and_b0_5  (\picorv32_core/sel43_b21/B5 , \picorv32_core/n525 [21], \picorv32_core/n664 );
  or \picorv32_core/sel43_b21/or_B2_B3  (\picorv32_core/sel43_b21/or_B2_B3_o , \picorv32_core/sel43_b21/B2 , \picorv32_core/sel43_b21/B3 );
  or \picorv32_core/sel43_b21/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b21/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b21/B0 , \picorv32_core/sel43_b21/or_B2_B3_o );
  or \picorv32_core/sel43_b21/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [21], \picorv32_core/sel43_b21/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b21/B5 );
  and \picorv32_core/sel43_b22/and_b0_0  (\picorv32_core/sel43_b22/B0 , \picorv32_core/n658 [22], \picorv32_core/n669 );
  and \picorv32_core/sel43_b22/and_b0_2  (\picorv32_core/sel43_b22/B2 , \picorv32_core/n567 [22], \picorv32_core/n667 );
  and \picorv32_core/sel43_b22/and_b0_3  (\picorv32_core/sel43_b22/B3 , \picorv32_core/n543 [22], \picorv32_core/n666 );
  and \picorv32_core/sel43_b22/and_b0_5  (\picorv32_core/sel43_b22/B5 , \picorv32_core/n525 [22], \picorv32_core/n664 );
  or \picorv32_core/sel43_b22/or_B2_B3  (\picorv32_core/sel43_b22/or_B2_B3_o , \picorv32_core/sel43_b22/B2 , \picorv32_core/sel43_b22/B3 );
  or \picorv32_core/sel43_b22/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b22/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b22/B0 , \picorv32_core/sel43_b22/or_B2_B3_o );
  or \picorv32_core/sel43_b22/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [22], \picorv32_core/sel43_b22/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b22/B5 );
  and \picorv32_core/sel43_b23/and_b0_0  (\picorv32_core/sel43_b23/B0 , \picorv32_core/n658 [23], \picorv32_core/n669 );
  and \picorv32_core/sel43_b23/and_b0_2  (\picorv32_core/sel43_b23/B2 , \picorv32_core/n567 [23], \picorv32_core/n667 );
  and \picorv32_core/sel43_b23/and_b0_3  (\picorv32_core/sel43_b23/B3 , \picorv32_core/n543 [23], \picorv32_core/n666 );
  and \picorv32_core/sel43_b23/and_b0_5  (\picorv32_core/sel43_b23/B5 , \picorv32_core/n525 [23], \picorv32_core/n664 );
  or \picorv32_core/sel43_b23/or_B2_B3  (\picorv32_core/sel43_b23/or_B2_B3_o , \picorv32_core/sel43_b23/B2 , \picorv32_core/sel43_b23/B3 );
  or \picorv32_core/sel43_b23/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b23/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b23/B0 , \picorv32_core/sel43_b23/or_B2_B3_o );
  or \picorv32_core/sel43_b23/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [23], \picorv32_core/sel43_b23/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b23/B5 );
  and \picorv32_core/sel43_b24/and_b0_0  (\picorv32_core/sel43_b24/B0 , \picorv32_core/n658 [24], \picorv32_core/n669 );
  and \picorv32_core/sel43_b24/and_b0_2  (\picorv32_core/sel43_b24/B2 , \picorv32_core/n567 [24], \picorv32_core/n667 );
  and \picorv32_core/sel43_b24/and_b0_3  (\picorv32_core/sel43_b24/B3 , \picorv32_core/n543 [24], \picorv32_core/n666 );
  and \picorv32_core/sel43_b24/and_b0_5  (\picorv32_core/sel43_b24/B5 , \picorv32_core/n525 [24], \picorv32_core/n664 );
  or \picorv32_core/sel43_b24/or_B2_B3  (\picorv32_core/sel43_b24/or_B2_B3_o , \picorv32_core/sel43_b24/B2 , \picorv32_core/sel43_b24/B3 );
  or \picorv32_core/sel43_b24/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b24/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b24/B0 , \picorv32_core/sel43_b24/or_B2_B3_o );
  or \picorv32_core/sel43_b24/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [24], \picorv32_core/sel43_b24/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b24/B5 );
  and \picorv32_core/sel43_b25/and_b0_0  (\picorv32_core/sel43_b25/B0 , \picorv32_core/n658 [25], \picorv32_core/n669 );
  and \picorv32_core/sel43_b25/and_b0_2  (\picorv32_core/sel43_b25/B2 , \picorv32_core/n567 [25], \picorv32_core/n667 );
  and \picorv32_core/sel43_b25/and_b0_3  (\picorv32_core/sel43_b25/B3 , \picorv32_core/n543 [25], \picorv32_core/n666 );
  and \picorv32_core/sel43_b25/and_b0_5  (\picorv32_core/sel43_b25/B5 , \picorv32_core/n525 [25], \picorv32_core/n664 );
  or \picorv32_core/sel43_b25/or_B2_B3  (\picorv32_core/sel43_b25/or_B2_B3_o , \picorv32_core/sel43_b25/B2 , \picorv32_core/sel43_b25/B3 );
  or \picorv32_core/sel43_b25/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b25/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b25/B0 , \picorv32_core/sel43_b25/or_B2_B3_o );
  or \picorv32_core/sel43_b25/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [25], \picorv32_core/sel43_b25/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b25/B5 );
  and \picorv32_core/sel43_b26/and_b0_0  (\picorv32_core/sel43_b26/B0 , \picorv32_core/n658 [26], \picorv32_core/n669 );
  and \picorv32_core/sel43_b26/and_b0_2  (\picorv32_core/sel43_b26/B2 , \picorv32_core/n567 [26], \picorv32_core/n667 );
  and \picorv32_core/sel43_b26/and_b0_3  (\picorv32_core/sel43_b26/B3 , \picorv32_core/n543 [26], \picorv32_core/n666 );
  and \picorv32_core/sel43_b26/and_b0_5  (\picorv32_core/sel43_b26/B5 , \picorv32_core/n525 [26], \picorv32_core/n664 );
  or \picorv32_core/sel43_b26/or_B2_B3  (\picorv32_core/sel43_b26/or_B2_B3_o , \picorv32_core/sel43_b26/B2 , \picorv32_core/sel43_b26/B3 );
  or \picorv32_core/sel43_b26/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b26/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b26/B0 , \picorv32_core/sel43_b26/or_B2_B3_o );
  or \picorv32_core/sel43_b26/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [26], \picorv32_core/sel43_b26/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b26/B5 );
  and \picorv32_core/sel43_b27/and_b0_0  (\picorv32_core/sel43_b27/B0 , \picorv32_core/n658 [27], \picorv32_core/n669 );
  and \picorv32_core/sel43_b27/and_b0_2  (\picorv32_core/sel43_b27/B2 , \picorv32_core/n567 [27], \picorv32_core/n667 );
  and \picorv32_core/sel43_b27/and_b0_3  (\picorv32_core/sel43_b27/B3 , \picorv32_core/n543 [27], \picorv32_core/n666 );
  and \picorv32_core/sel43_b27/and_b0_5  (\picorv32_core/sel43_b27/B5 , \picorv32_core/n525 [27], \picorv32_core/n664 );
  or \picorv32_core/sel43_b27/or_B2_B3  (\picorv32_core/sel43_b27/or_B2_B3_o , \picorv32_core/sel43_b27/B2 , \picorv32_core/sel43_b27/B3 );
  or \picorv32_core/sel43_b27/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b27/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b27/B0 , \picorv32_core/sel43_b27/or_B2_B3_o );
  or \picorv32_core/sel43_b27/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [27], \picorv32_core/sel43_b27/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b27/B5 );
  and \picorv32_core/sel43_b28/and_b0_0  (\picorv32_core/sel43_b28/B0 , \picorv32_core/n658 [28], \picorv32_core/n669 );
  and \picorv32_core/sel43_b28/and_b0_2  (\picorv32_core/sel43_b28/B2 , \picorv32_core/n567 [28], \picorv32_core/n667 );
  and \picorv32_core/sel43_b28/and_b0_3  (\picorv32_core/sel43_b28/B3 , \picorv32_core/n543 [28], \picorv32_core/n666 );
  and \picorv32_core/sel43_b28/and_b0_5  (\picorv32_core/sel43_b28/B5 , \picorv32_core/n525 [28], \picorv32_core/n664 );
  or \picorv32_core/sel43_b28/or_B2_B3  (\picorv32_core/sel43_b28/or_B2_B3_o , \picorv32_core/sel43_b28/B2 , \picorv32_core/sel43_b28/B3 );
  or \picorv32_core/sel43_b28/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b28/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b28/B0 , \picorv32_core/sel43_b28/or_B2_B3_o );
  or \picorv32_core/sel43_b28/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [28], \picorv32_core/sel43_b28/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b28/B5 );
  and \picorv32_core/sel43_b29/and_b0_0  (\picorv32_core/sel43_b29/B0 , \picorv32_core/n658 [29], \picorv32_core/n669 );
  and \picorv32_core/sel43_b29/and_b0_2  (\picorv32_core/sel43_b29/B2 , \picorv32_core/n567 [29], \picorv32_core/n667 );
  and \picorv32_core/sel43_b29/and_b0_3  (\picorv32_core/sel43_b29/B3 , \picorv32_core/n543 [29], \picorv32_core/n666 );
  and \picorv32_core/sel43_b29/and_b0_5  (\picorv32_core/sel43_b29/B5 , \picorv32_core/n525 [29], \picorv32_core/n664 );
  or \picorv32_core/sel43_b29/or_B2_B3  (\picorv32_core/sel43_b29/or_B2_B3_o , \picorv32_core/sel43_b29/B2 , \picorv32_core/sel43_b29/B3 );
  or \picorv32_core/sel43_b29/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b29/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b29/B0 , \picorv32_core/sel43_b29/or_B2_B3_o );
  or \picorv32_core/sel43_b29/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [29], \picorv32_core/sel43_b29/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b29/B5 );
  and \picorv32_core/sel43_b3/and_b0_0  (\picorv32_core/sel43_b3/B0 , \picorv32_core/n658 [3], \picorv32_core/n669 );
  and \picorv32_core/sel43_b3/and_b0_2  (\picorv32_core/sel43_b3/B2 , \picorv32_core/n567 [3], \picorv32_core/n667 );
  and \picorv32_core/sel43_b3/and_b0_3  (\picorv32_core/sel43_b3/B3 , \picorv32_core/n543 [3], \picorv32_core/n666 );
  and \picorv32_core/sel43_b3/and_b0_5  (\picorv32_core/sel43_b3/B5 , \picorv32_core/n525 [3], \picorv32_core/n664 );
  or \picorv32_core/sel43_b3/or_B2_B3  (\picorv32_core/sel43_b3/or_B2_B3_o , \picorv32_core/sel43_b3/B2 , \picorv32_core/sel43_b3/B3 );
  or \picorv32_core/sel43_b3/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b3/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b3/B0 , \picorv32_core/sel43_b3/or_B2_B3_o );
  or \picorv32_core/sel43_b3/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [3], \picorv32_core/sel43_b3/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b3/B5 );
  and \picorv32_core/sel43_b30/and_b0_0  (\picorv32_core/sel43_b30/B0 , \picorv32_core/n658 [30], \picorv32_core/n669 );
  and \picorv32_core/sel43_b30/and_b0_2  (\picorv32_core/sel43_b30/B2 , \picorv32_core/n567 [30], \picorv32_core/n667 );
  and \picorv32_core/sel43_b30/and_b0_3  (\picorv32_core/sel43_b30/B3 , \picorv32_core/n543 [30], \picorv32_core/n666 );
  and \picorv32_core/sel43_b30/and_b0_5  (\picorv32_core/sel43_b30/B5 , \picorv32_core/n525 [30], \picorv32_core/n664 );
  or \picorv32_core/sel43_b30/or_B2_B3  (\picorv32_core/sel43_b30/or_B2_B3_o , \picorv32_core/sel43_b30/B2 , \picorv32_core/sel43_b30/B3 );
  or \picorv32_core/sel43_b30/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b30/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b30/B0 , \picorv32_core/sel43_b30/or_B2_B3_o );
  or \picorv32_core/sel43_b30/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [30], \picorv32_core/sel43_b30/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b30/B5 );
  and \picorv32_core/sel43_b31/and_b0_0  (\picorv32_core/sel43_b31/B0 , \picorv32_core/n658 [31], \picorv32_core/n669 );
  and \picorv32_core/sel43_b31/and_b0_2  (\picorv32_core/sel43_b31/B2 , \picorv32_core/n567 [31], \picorv32_core/n667 );
  and \picorv32_core/sel43_b31/and_b0_3  (\picorv32_core/sel43_b31/B3 , \picorv32_core/n543 [31], \picorv32_core/n666 );
  and \picorv32_core/sel43_b31/and_b0_5  (\picorv32_core/sel43_b31/B5 , \picorv32_core/n525 [31], \picorv32_core/n664 );
  or \picorv32_core/sel43_b31/or_B2_B3  (\picorv32_core/sel43_b31/or_B2_B3_o , \picorv32_core/sel43_b31/B2 , \picorv32_core/sel43_b31/B3 );
  or \picorv32_core/sel43_b31/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b31/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b31/B0 , \picorv32_core/sel43_b31/or_B2_B3_o );
  or \picorv32_core/sel43_b31/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [31], \picorv32_core/sel43_b31/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b31/B5 );
  and \picorv32_core/sel43_b4/and_b0_0  (\picorv32_core/sel43_b4/B0 , \picorv32_core/n658 [4], \picorv32_core/n669 );
  and \picorv32_core/sel43_b4/and_b0_2  (\picorv32_core/sel43_b4/B2 , \picorv32_core/n567 [4], \picorv32_core/n667 );
  and \picorv32_core/sel43_b4/and_b0_3  (\picorv32_core/sel43_b4/B3 , \picorv32_core/n543 [4], \picorv32_core/n666 );
  and \picorv32_core/sel43_b4/and_b0_5  (\picorv32_core/sel43_b4/B5 , \picorv32_core/n525 [4], \picorv32_core/n664 );
  or \picorv32_core/sel43_b4/or_B2_B3  (\picorv32_core/sel43_b4/or_B2_B3_o , \picorv32_core/sel43_b4/B2 , \picorv32_core/sel43_b4/B3 );
  or \picorv32_core/sel43_b4/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b4/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b4/B0 , \picorv32_core/sel43_b4/or_B2_B3_o );
  or \picorv32_core/sel43_b4/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [4], \picorv32_core/sel43_b4/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b4/B5 );
  and \picorv32_core/sel43_b5/and_b0_0  (\picorv32_core/sel43_b5/B0 , \picorv32_core/n658 [5], \picorv32_core/n669 );
  and \picorv32_core/sel43_b5/and_b0_2  (\picorv32_core/sel43_b5/B2 , \picorv32_core/n567 [5], \picorv32_core/n667 );
  and \picorv32_core/sel43_b5/and_b0_3  (\picorv32_core/sel43_b5/B3 , \picorv32_core/n543 [5], \picorv32_core/n666 );
  and \picorv32_core/sel43_b5/and_b0_5  (\picorv32_core/sel43_b5/B5 , \picorv32_core/n525 [5], \picorv32_core/n664 );
  or \picorv32_core/sel43_b5/or_B2_B3  (\picorv32_core/sel43_b5/or_B2_B3_o , \picorv32_core/sel43_b5/B2 , \picorv32_core/sel43_b5/B3 );
  or \picorv32_core/sel43_b5/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b5/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b5/B0 , \picorv32_core/sel43_b5/or_B2_B3_o );
  or \picorv32_core/sel43_b5/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [5], \picorv32_core/sel43_b5/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b5/B5 );
  and \picorv32_core/sel43_b6/and_b0_0  (\picorv32_core/sel43_b6/B0 , \picorv32_core/n658 [6], \picorv32_core/n669 );
  and \picorv32_core/sel43_b6/and_b0_2  (\picorv32_core/sel43_b6/B2 , \picorv32_core/n567 [6], \picorv32_core/n667 );
  and \picorv32_core/sel43_b6/and_b0_3  (\picorv32_core/sel43_b6/B3 , \picorv32_core/n543 [6], \picorv32_core/n666 );
  and \picorv32_core/sel43_b6/and_b0_5  (\picorv32_core/sel43_b6/B5 , \picorv32_core/n525 [6], \picorv32_core/n664 );
  or \picorv32_core/sel43_b6/or_B2_B3  (\picorv32_core/sel43_b6/or_B2_B3_o , \picorv32_core/sel43_b6/B2 , \picorv32_core/sel43_b6/B3 );
  or \picorv32_core/sel43_b6/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b6/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b6/B0 , \picorv32_core/sel43_b6/or_B2_B3_o );
  or \picorv32_core/sel43_b6/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [6], \picorv32_core/sel43_b6/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b6/B5 );
  and \picorv32_core/sel43_b7/and_b0_0  (\picorv32_core/sel43_b7/B0 , \picorv32_core/n658 [7], \picorv32_core/n669 );
  and \picorv32_core/sel43_b7/and_b0_2  (\picorv32_core/sel43_b7/B2 , \picorv32_core/n567 [7], \picorv32_core/n667 );
  and \picorv32_core/sel43_b7/and_b0_3  (\picorv32_core/sel43_b7/B3 , \picorv32_core/n543 [7], \picorv32_core/n666 );
  and \picorv32_core/sel43_b7/and_b0_5  (\picorv32_core/sel43_b7/B5 , \picorv32_core/n525 [7], \picorv32_core/n664 );
  or \picorv32_core/sel43_b7/or_B2_B3  (\picorv32_core/sel43_b7/or_B2_B3_o , \picorv32_core/sel43_b7/B2 , \picorv32_core/sel43_b7/B3 );
  or \picorv32_core/sel43_b7/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b7/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b7/B0 , \picorv32_core/sel43_b7/or_B2_B3_o );
  or \picorv32_core/sel43_b7/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [7], \picorv32_core/sel43_b7/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b7/B5 );
  and \picorv32_core/sel43_b8/and_b0_0  (\picorv32_core/sel43_b8/B0 , \picorv32_core/n658 [8], \picorv32_core/n669 );
  and \picorv32_core/sel43_b8/and_b0_2  (\picorv32_core/sel43_b8/B2 , \picorv32_core/n567 [8], \picorv32_core/n667 );
  and \picorv32_core/sel43_b8/and_b0_3  (\picorv32_core/sel43_b8/B3 , \picorv32_core/n543 [8], \picorv32_core/n666 );
  and \picorv32_core/sel43_b8/and_b0_5  (\picorv32_core/sel43_b8/B5 , \picorv32_core/n525 [8], \picorv32_core/n664 );
  or \picorv32_core/sel43_b8/or_B2_B3  (\picorv32_core/sel43_b8/or_B2_B3_o , \picorv32_core/sel43_b8/B2 , \picorv32_core/sel43_b8/B3 );
  or \picorv32_core/sel43_b8/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b8/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b8/B0 , \picorv32_core/sel43_b8/or_B2_B3_o );
  or \picorv32_core/sel43_b8/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [8], \picorv32_core/sel43_b8/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b8/B5 );
  and \picorv32_core/sel43_b9/and_b0_0  (\picorv32_core/sel43_b9/B0 , \picorv32_core/n658 [9], \picorv32_core/n669 );
  and \picorv32_core/sel43_b9/and_b0_2  (\picorv32_core/sel43_b9/B2 , \picorv32_core/n567 [9], \picorv32_core/n667 );
  and \picorv32_core/sel43_b9/and_b0_3  (\picorv32_core/sel43_b9/B3 , \picorv32_core/n543 [9], \picorv32_core/n666 );
  and \picorv32_core/sel43_b9/and_b0_5  (\picorv32_core/sel43_b9/B5 , \picorv32_core/n525 [9], \picorv32_core/n664 );
  or \picorv32_core/sel43_b9/or_B2_B3  (\picorv32_core/sel43_b9/or_B2_B3_o , \picorv32_core/sel43_b9/B2 , \picorv32_core/sel43_b9/B3 );
  or \picorv32_core/sel43_b9/or_or_B0_B1_o_or_B2_  (\picorv32_core/sel43_b9/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b9/B0 , \picorv32_core/sel43_b9/or_B2_B3_o );
  or \picorv32_core/sel43_b9/or_or_or_B0_B1_o_or_  (\picorv32_core/n695 [9], \picorv32_core/sel43_b9/or_or_B0_B1_o_or_B2__o , \picorv32_core/sel43_b9/B5 );
  and \picorv32_core/sel44_b0/and_b0_2  (\picorv32_core/sel44_b0/B2 , \picorv32_core/n571 [0], \picorv32_core/n667 );
  and \picorv32_core/sel44_b0/and_b0_5  (\picorv32_core/sel44_b0/B5 , \picorv32_core/n532 [0], \picorv32_core/n664 );
  or \picorv32_core/sel44_b0/or_B4_B5  (\picorv32_core/sel44_b0/or_B4_B5_o , \picorv32_core/sel42_b0/B4 , \picorv32_core/sel44_b0/B5 );
  or \picorv32_core/sel44_b0/or_or_or_B0_B1_o_or_  (\picorv32_core/n696 [0], \picorv32_core/sel44_b0/B2 , \picorv32_core/sel44_b0/or_B4_B5_o );
  and \picorv32_core/sel44_b1/and_b0_2  (\picorv32_core/sel44_b1/B2 , \picorv32_core/n571 [1], \picorv32_core/n667 );
  and \picorv32_core/sel44_b1/and_b0_5  (\picorv32_core/sel44_b1/B5 , \picorv32_core/n532 [1], \picorv32_core/n664 );
  or \picorv32_core/sel44_b1/or_B4_B5  (\picorv32_core/sel44_b1/or_B4_B5_o , \picorv32_core/sel42_b1/B4 , \picorv32_core/sel44_b1/B5 );
  or \picorv32_core/sel44_b1/or_or_or_B0_B1_o_or_  (\picorv32_core/n696 [1], \picorv32_core/sel44_b1/B2 , \picorv32_core/sel44_b1/or_B4_B5_o );
  and \picorv32_core/sel44_b2/and_b0_2  (\picorv32_core/sel44_b2/B2 , \picorv32_core/n571 [2], \picorv32_core/n667 );
  and \picorv32_core/sel44_b2/and_b0_5  (\picorv32_core/sel44_b2/B5 , \picorv32_core/n532 [2], \picorv32_core/n664 );
  or \picorv32_core/sel44_b2/or_B4_B5  (\picorv32_core/sel44_b2/or_B4_B5_o , \picorv32_core/sel42_b2/B4 , \picorv32_core/sel44_b2/B5 );
  or \picorv32_core/sel44_b2/or_or_or_B0_B1_o_or_  (\picorv32_core/n696 [2], \picorv32_core/sel44_b2/B2 , \picorv32_core/sel44_b2/or_B4_B5_o );
  and \picorv32_core/sel44_b3/and_b0_2  (\picorv32_core/sel44_b3/B2 , \picorv32_core/n571 [3], \picorv32_core/n667 );
  and \picorv32_core/sel44_b3/and_b0_5  (\picorv32_core/sel44_b3/B5 , \picorv32_core/n532 [3], \picorv32_core/n664 );
  or \picorv32_core/sel44_b3/or_B4_B5  (\picorv32_core/sel44_b3/or_B4_B5_o , \picorv32_core/sel42_b3/B4 , \picorv32_core/sel44_b3/B5 );
  or \picorv32_core/sel44_b3/or_or_or_B0_B1_o_or_  (\picorv32_core/n696 [3], \picorv32_core/sel44_b3/B2 , \picorv32_core/sel44_b3/or_B4_B5_o );
  and \picorv32_core/sel44_b4/and_b0_2  (\picorv32_core/sel44_b4/B2 , \picorv32_core/n571 [4], \picorv32_core/n667 );
  and \picorv32_core/sel44_b4/and_b0_5  (\picorv32_core/sel44_b4/B5 , \picorv32_core/n532 [4], \picorv32_core/n664 );
  or \picorv32_core/sel44_b4/or_B4_B5  (\picorv32_core/sel44_b4/or_B4_B5_o , \picorv32_core/sel42_b4/B4 , \picorv32_core/sel44_b4/B5 );
  or \picorv32_core/sel44_b4/or_or_or_B0_B1_o_or_  (\picorv32_core/n696 [4], \picorv32_core/sel44_b4/B2 , \picorv32_core/sel44_b4/or_B4_B5_o );
  and \picorv32_core/sel45/and_b0_0  (\picorv32_core/sel45/B0 , \picorv32_core/n659 , \picorv32_core/n669 );
  and \picorv32_core/sel45/and_b0_1  (\picorv32_core/sel45/B1 , \picorv32_core/n659 , \picorv32_core/n668 );
  and \picorv32_core/sel45/and_b0_2  (\picorv32_core/sel45/B2 , \picorv32_core/n550 , \picorv32_core/n666 );
  and \picorv32_core/sel45/and_b0_3  (\picorv32_core/sel45/B3 , \picorv32_core/n170 , \picorv32_core/n697 );
  or \picorv32_core/sel45/or_B0_B1  (\picorv32_core/sel45/or_B0_B1_o , \picorv32_core/sel45/B0 , \picorv32_core/sel45/B1 );
  or \picorv32_core/sel45/or_B2_B3  (\picorv32_core/sel45/or_B2_B3_o , \picorv32_core/sel45/B2 , \picorv32_core/sel45/B3 );
  or \picorv32_core/sel45/or_or_B0_B1_o_or_B2_  (\picorv32_core/n698 , \picorv32_core/sel45/or_B0_B1_o , \picorv32_core/sel45/or_B2_B3_o );
  and \picorv32_core/sel46_sel_is_2  (\picorv32_core/sel46_sel_is_2_o , \picorv32_core/n701_neg , \picorv32_core/n597 );
  and \picorv32_core/sel4_b0/and_b0_0  (\picorv32_core/sel4_b0/B0 , \picorv32_core/n42 [12], \picorv32_core/n100 );
  and \picorv32_core/sel4_b0/and_b0_1  (\picorv32_core/sel4_b0/B1 , \picorv32_core/n95 [0], \picorv32_core/n98 );
  or \picorv32_core/sel4_b0/or_B0_B1  (\picorv32_core/sel4_b0/or_B0_B1_o , \picorv32_core/sel4_b0/B0 , \picorv32_core/sel4_b0/B1 );
  or \picorv32_core/sel4_b0/or_or_B0_B1_o_or_B2_  (\picorv32_core/n105 [0], \picorv32_core/sel4_b0/or_B0_B1_o , \picorv32_core/n96 );
  and \picorv32_core/sel4_b1/and_b0_0  (\picorv32_core/sel4_b1/B0 , \picorv32_core/n42 [13], \picorv32_core/n100 );
  and \picorv32_core/sel4_b1/and_b0_1  (\picorv32_core/sel4_b1/B1 , \picorv32_core/n95 [1], \picorv32_core/n98 );
  or \picorv32_core/sel4_b1/or_B0_B1  (\picorv32_core/sel4_b1/or_B0_B1_o , \picorv32_core/sel4_b1/B0 , \picorv32_core/sel4_b1/B1 );
  or \picorv32_core/sel4_b1/or_or_B0_B1_o_or_B2_  (\picorv32_core/n105 [1], \picorv32_core/sel4_b1/or_B0_B1_o , \picorv32_core/n104 );
  and \picorv32_core/sel4_b2/and_b0_0  (\picorv32_core/sel4_b2/B0 , \picorv32_core/n42 [25], \picorv32_core/n100 );
  and \picorv32_core/sel4_b2/and_b0_1  (\picorv32_core/sel4_b2/B1 , \picorv32_core/n95 [2], \picorv32_core/n98 );
  and \picorv32_core/sel4_b2/and_b0_2  (\picorv32_core/sel4_b2/B2 , \picorv32_core/mem_rdata_latched [12], \picorv32_core/n104 );
  or \picorv32_core/sel4_b2/or_B0_B1  (\picorv32_core/sel4_b2/or_B0_B1_o , \picorv32_core/sel4_b2/B0 , \picorv32_core/sel4_b2/B1 );
  or \picorv32_core/sel4_b2/or_or_B0_B1_o_or_B2_  (\picorv32_core/n105 [2], \picorv32_core/sel4_b2/or_B0_B1_o , \picorv32_core/sel4_b2/B2 );
  and \picorv32_core/sel5_b0/and_b0_0  (\picorv32_core/sel5_b0/B0 , \picorv32_core/n91 [0], \picorv32_core/n98 );
  and \picorv32_core/sel5_b0/and_b0_2  (\picorv32_core/sel5_b0/B2 , \picorv32_core/n42 [20], \picorv32_core/n106 );
  or \picorv32_core/sel5_b0/or_B0_or_B1_B2_o  (\picorv32_core/n107 [0], \picorv32_core/sel5_b0/B0 , \picorv32_core/sel5_b0/B2 );
  and \picorv32_core/sel5_b1/and_b0_0  (\picorv32_core/sel5_b1/B0 , \picorv32_core/n91 [1], \picorv32_core/n98 );
  and \picorv32_core/sel5_b1/and_b0_2  (\picorv32_core/sel5_b1/B2 , \picorv32_core/n42 [21], \picorv32_core/n106 );
  or \picorv32_core/sel5_b1/or_B0_or_B1_B2_o  (\picorv32_core/n107 [1], \picorv32_core/sel5_b1/B0 , \picorv32_core/sel5_b1/B2 );
  and \picorv32_core/sel5_b2/and_b0_0  (\picorv32_core/sel5_b2/B0 , \picorv32_core/n91 [2], \picorv32_core/n98 );
  and \picorv32_core/sel5_b2/and_b0_1  (\picorv32_core/sel5_b2/B1 , \picorv32_core/mem_rdata_latched [4], \picorv32_core/n97 );
  and \picorv32_core/sel5_b2/and_b0_2  (\picorv32_core/sel5_b2/B2 , \picorv32_core/n42 [22], \picorv32_core/n106 );
  or \picorv32_core/sel5_b2/or_B0_or_B1_B2_o  (\picorv32_core/n107 [2], \picorv32_core/sel5_b2/B0 , \picorv32_core/sel5_b2/or_B1_B2_o );
  or \picorv32_core/sel5_b2/or_B1_B2  (\picorv32_core/sel5_b2/or_B1_B2_o , \picorv32_core/sel5_b2/B1 , \picorv32_core/sel5_b2/B2 );
  and \picorv32_core/sel5_b3/and_b0_0  (\picorv32_core/sel5_b3/B0 , \picorv32_core/n91 [3], \picorv32_core/n98 );
  and \picorv32_core/sel5_b3/and_b0_1  (\picorv32_core/sel5_b3/B1 , \picorv32_core/mem_rdata_latched [5], \picorv32_core/n97 );
  and \picorv32_core/sel5_b3/and_b0_2  (\picorv32_core/sel5_b3/B2 , \picorv32_core/n42 [23], \picorv32_core/n106 );
  or \picorv32_core/sel5_b3/or_B0_or_B1_B2_o  (\picorv32_core/n107 [3], \picorv32_core/sel5_b3/B0 , \picorv32_core/sel5_b3/or_B1_B2_o );
  or \picorv32_core/sel5_b3/or_B1_B2  (\picorv32_core/sel5_b3/or_B1_B2_o , \picorv32_core/sel5_b3/B1 , \picorv32_core/sel5_b3/B2 );
  and \picorv32_core/sel5_b4/and_b0_0  (\picorv32_core/sel5_b4/B0 , \picorv32_core/n91 [4], \picorv32_core/n98 );
  and \picorv32_core/sel5_b4/and_b0_1  (\picorv32_core/sel5_b4/B1 , \picorv32_core/mem_rdata_latched [6], \picorv32_core/n97 );
  and \picorv32_core/sel5_b4/and_b0_2  (\picorv32_core/sel5_b4/B2 , \picorv32_core/n42 [24], \picorv32_core/n106 );
  or \picorv32_core/sel5_b4/or_B0_or_B1_B2_o  (\picorv32_core/n107 [4], \picorv32_core/sel5_b4/B0 , \picorv32_core/sel5_b4/or_B1_B2_o );
  or \picorv32_core/sel5_b4/or_B1_B2  (\picorv32_core/sel5_b4/or_B1_B2_o , \picorv32_core/sel5_b4/B1 , \picorv32_core/sel5_b4/B2 );
  and \picorv32_core/sel6_b0/and_b0_0  (\picorv32_core/sel6_b0/B0 , \picorv32_core/n42 [13], \picorv32_core/n44 );
  or \picorv32_core/sel6_b0/or_B0_or_B1_B2_o  (\picorv32_core/n47 [0], \picorv32_core/sel6_b0/B0 , \picorv32_core/n104 );
  and \picorv32_core/sel6_b1/and_b0_0  (\picorv32_core/sel6_b1/B0 , \picorv32_core/n42 [26], \picorv32_core/n44 );
  and \picorv32_core/sel6_b1/and_b0_1  (\picorv32_core/sel6_b1/B1 , \picorv32_core/mem_rdata_latched [5], \picorv32_core/n104 );
  and \picorv32_core/sel6_b1/and_b0_2  (\picorv32_core/sel6_b1/B2 , \picorv32_core/mem_rdata_latched [7], \picorv32_core/n96 );
  or \picorv32_core/sel6_b1/or_B0_or_B1_B2_o  (\picorv32_core/n47 [1], \picorv32_core/sel6_b1/B0 , \picorv32_core/sel6_b1/or_B1_B2_o );
  or \picorv32_core/sel6_b1/or_B1_B2  (\picorv32_core/sel6_b1/or_B1_B2_o , \picorv32_core/sel6_b1/B1 , \picorv32_core/sel6_b1/B2 );
  and \picorv32_core/sel6_b2/and_b0_0  (\picorv32_core/sel6_b2/B0 , \picorv32_core/n42 [27], \picorv32_core/n44 );
  and \picorv32_core/sel6_b2/and_b0_2  (\picorv32_core/sel6_b2/B2 , \picorv32_core/mem_rdata_latched [8], \picorv32_core/n96 );
  or \picorv32_core/sel6_b2/or_B0_or_B1_B2_o  (\picorv32_core/n47 [2], \picorv32_core/sel6_b2/B0 , \picorv32_core/sel6_b2/B2 );
  and \picorv32_core/sel6_b3/and_b0_0  (\picorv32_core/sel6_b3/B0 , \picorv32_core/n42 [28], \picorv32_core/n44 );
  and \picorv32_core/sel6_b3/and_b0_2  (\picorv32_core/sel6_b3/B2 , \picorv32_core/mem_rdata_latched [9], \picorv32_core/n96 );
  or \picorv32_core/sel6_b3/or_B0_or_B1_B2_o  (\picorv32_core/n47 [3], \picorv32_core/sel6_b3/B0 , \picorv32_core/sel6_b3/B2 );
  and \picorv32_core/sel6_b4/and_b0_0  (\picorv32_core/sel6_b4/B0 , \picorv32_core/n42 [29], \picorv32_core/n44 );
  and \picorv32_core/sel6_b4/and_b0_2  (\picorv32_core/sel6_b4/B2 , \picorv32_core/mem_rdata_latched [10], \picorv32_core/n96 );
  or \picorv32_core/sel6_b4/or_B0_or_B1_B2_o  (\picorv32_core/n47 [4], \picorv32_core/sel6_b4/B0 , \picorv32_core/sel6_b4/B2 );
  and \picorv32_core/sel7/and_b0_1  (\picorv32_core/sel7/B1 , \picorv32_core/mem_rdata_latched [8], \picorv32_core/n104 );
  or \picorv32_core/sel7/or_B1_B2  (\picorv32_core/sel7/or_B1_B2_o , \picorv32_core/sel7/B1 , \picorv32_core/n96 );
  binary_mux_s3_w1 \picorv32_core/sel8_b0  (
    .i0(\picorv32_core/mem_rdata_latched [7]),
    .i1(1'b0),
    .i2(\picorv32_core/mem_rdata_latched [7]),
    .i3(1'b0),
    .i4(\picorv32_core/n225 [0]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n229 [0]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel8_b1  (
    .i0(\picorv32_core/mem_rdata_latched [8]),
    .i1(1'b0),
    .i2(\picorv32_core/mem_rdata_latched [8]),
    .i3(1'b0),
    .i4(\picorv32_core/n225 [1]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n229 [1]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel8_b2  (
    .i0(\picorv32_core/mem_rdata_latched [9]),
    .i1(1'b0),
    .i2(\picorv32_core/mem_rdata_latched [9]),
    .i3(1'b0),
    .i4(\picorv32_core/n225 [2]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n229 [2]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel8_b3  (
    .i0(\picorv32_core/mem_rdata_latched [10]),
    .i1(1'b0),
    .i2(\picorv32_core/mem_rdata_latched [10]),
    .i3(1'b0),
    .i4(\picorv32_core/n225 [3]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n229 [3]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel8_b4  (
    .i0(\picorv32_core/mem_rdata_latched [11]),
    .i1(1'b0),
    .i2(\picorv32_core/mem_rdata_latched [11]),
    .i3(1'b0),
    .i4(\picorv32_core/n225 [4]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n229 [4]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel9_b0  (
    .i0(\picorv32_core/mem_rdata_latched [7]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\picorv32_core/n226 [0]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n230 [0]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel9_b1  (
    .i0(\picorv32_core/mem_rdata_latched [8]),
    .i1(1'b0),
    .i2(1'b1),
    .i3(1'b0),
    .i4(\picorv32_core/n226 [1]),
    .i5(1'b0),
    .i6(1'b1),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n230 [1]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel9_b2  (
    .i0(\picorv32_core/mem_rdata_latched [9]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\picorv32_core/n226 [2]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n230 [2]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel9_b3  (
    .i0(\picorv32_core/mem_rdata_latched [10]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\picorv32_core/n226 [3]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n230 [3]));  // ../src/picorv32.v(987)
  binary_mux_s3_w1 \picorv32_core/sel9_b4  (
    .i0(\picorv32_core/mem_rdata_latched [11]),
    .i1(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\picorv32_core/n226 [4]),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\picorv32_core/mem_rdata_latched [15:13]),
    .o(\picorv32_core/n230 [4]));  // ../src/picorv32.v(987)
  add_pu32_mu32_o32 \picorv32_core/sub0  (
    .i0({\picorv32_core/pcpi_rs1$31$ ,\picorv32_core/pcpi_rs1$30$ ,\picorv32_core/pcpi_rs1$29$ ,\picorv32_core/pcpi_rs1$28$ ,\picorv32_core/pcpi_rs1$27$ ,\picorv32_core/pcpi_rs1$26$ ,\picorv32_core/pcpi_rs1$25$ ,\picorv32_core/pcpi_rs1$24$ ,\picorv32_core/pcpi_rs1$23$ ,\picorv32_core/pcpi_rs1$22$ ,\picorv32_core/pcpi_rs1$21$ ,\picorv32_core/pcpi_rs1$20$ ,\picorv32_core/pcpi_rs1$19$ ,\picorv32_core/pcpi_rs1$18$ ,\picorv32_core/pcpi_rs1$17$ ,\picorv32_core/pcpi_rs1$16$ ,\picorv32_core/pcpi_rs1$15$ ,\picorv32_core/pcpi_rs1$14$ ,\picorv32_core/pcpi_rs1$13$ ,\picorv32_core/pcpi_rs1$12$ ,\picorv32_core/pcpi_rs1$11$ ,\picorv32_core/pcpi_rs1$10$ ,\picorv32_core/pcpi_rs1$9$ ,\picorv32_core/pcpi_rs1$8$ ,\picorv32_core/pcpi_rs1$7$ ,\picorv32_core/pcpi_rs1$6$ ,\picorv32_core/pcpi_rs1$5$ ,\picorv32_core/pcpi_rs1$4$ ,\picorv32_core/pcpi_rs1$3$ ,\picorv32_core/pcpi_rs1$2$ ,\picorv32_core/pcpi_rs1$1$ ,\picorv32_core/pcpi_rs1$0$ }),
    .i1({\picorv32_core/pcpi_rs2$31$ ,\picorv32_core/pcpi_rs2$30$ ,\picorv32_core/pcpi_rs2$29$ ,\picorv32_core/pcpi_rs2$28$ ,\picorv32_core/pcpi_rs2$27$ ,\picorv32_core/pcpi_rs2$26$ ,\picorv32_core/pcpi_rs2$25$ ,\picorv32_core/pcpi_rs2$24$ ,\picorv32_core/pcpi_rs2$23$ ,\picorv32_core/pcpi_rs2$22$ ,\picorv32_core/pcpi_rs2$21$ ,\picorv32_core/pcpi_rs2$20$ ,\picorv32_core/pcpi_rs2$19$ ,\picorv32_core/pcpi_rs2$18$ ,\picorv32_core/pcpi_rs2$17$ ,\picorv32_core/pcpi_rs2$16$ ,\picorv32_core/pcpi_rs2$15$ ,\picorv32_core/pcpi_rs2$14$ ,\picorv32_core/pcpi_rs2$13$ ,\picorv32_core/pcpi_rs2$12$ ,\picorv32_core/pcpi_rs2$11$ ,\picorv32_core/pcpi_rs2$10$ ,\picorv32_core/pcpi_rs2$9$ ,\picorv32_core/pcpi_rs2$8$ ,mem_la_wdata[7:0]}),
    .o(\picorv32_core/n433 ));  // ../src/picorv32.v(1193)
  add_pu5_mu5_o5 \picorv32_core/sub1  (
    .i0(\picorv32_core/reg_sh ),
    .i1(5'b00100),
    .o(\picorv32_core/n559 [4:0]));  // ../src/picorv32.v(1780)
  add_pu5_mu5_o5 \picorv32_core/sub2  (
    .i0(\picorv32_core/reg_sh ),
    .i1(5'b00001),
    .o(\picorv32_core/n564 [4:0]));  // ../src/picorv32.v(1788)
  reg_sr_as_w1 \picorv32_core/trap_reg  (
    .clk(clk),
    .d(\picorv32_core/n662 ),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(trap));  // ../src/picorv32.v(1906)
  and \picorv32_core/u10  (\picorv32_core/mem_la_firstword_xfer , \picorv32_core/mem_xfer , \picorv32_core/mem_la_firstword );  // ../src/picorv32.v(327)
  and \picorv32_core/u100  (\picorv32_core/n87 , \picorv32_core/n86 , \picorv32_core/n73 );  // ../src/picorv32.v(491)
  and \picorv32_core/u101  (\picorv32_core/n443 [6], \picorv32_core/pcpi_rs1$6$ , mem_la_wdata[6]);  // ../src/picorv32.v(1232)
  and \picorv32_core/u102  (\picorv32_core/n443 [7], \picorv32_core/pcpi_rs1$7$ , mem_la_wdata[7]);  // ../src/picorv32.v(1232)
  and \picorv32_core/u103  (\picorv32_core/n443 [8], \picorv32_core/pcpi_rs1$8$ , \picorv32_core/pcpi_rs2$8$ );  // ../src/picorv32.v(1232)
  or \picorv32_core/u104  (\picorv32_core/n595 , \picorv32_core/n669 , \picorv32_core/n594 );  // ../src/picorv32.v(1851)
  or \picorv32_core/u105  (\picorv32_core/n37 , \picorv32_core/n664 , \picorv32_core/n662 );  // ../src/picorv32.v(1851)
  or \picorv32_core/u106  (\picorv32_core/n746 , \picorv32_core/n665 , \picorv32_core/n37 );  // ../src/picorv32.v(1851)
  or \picorv32_core/u107  (\picorv32_core/n678 , \picorv32_core/n595 , \picorv32_core/n746 );  // ../src/picorv32.v(1851)
  and \picorv32_core/u108  (\picorv32_core/n443 [9], \picorv32_core/pcpi_rs1$9$ , \picorv32_core/pcpi_rs2$9$ );  // ../src/picorv32.v(1232)
  not \picorv32_core/u109  (\picorv32_core/n523 , \picorv32_core/n647 );  // ../src/picorv32.v(1694)
  and \picorv32_core/u11  (\picorv32_core/n4 , \picorv32_core/mem_la_firstword , \picorv32_core/prefetched_high_word );  // ../src/picorv32.v(336)
  not \picorv32_core/u110  (\picorv32_core/n520 , \picorv32_core/n646 );  // ../src/picorv32.v(1690)
  and \picorv32_core/u113  (\picorv32_core/n92 , \picorv32_core/n84 , \picorv32_core/n79 );  // ../src/picorv32.v(495)
  and \picorv32_core/u114  (\picorv32_core/n443 [10], \picorv32_core/pcpi_rs1$10$ , \picorv32_core/pcpi_rs2$10$ );  // ../src/picorv32.v(1232)
  and \picorv32_core/u115  (\picorv32_core/n443 [11], \picorv32_core/pcpi_rs1$11$ , \picorv32_core/pcpi_rs2$11$ );  // ../src/picorv32.v(1232)
  and \picorv32_core/u116  (\picorv32_core/n443 [12], \picorv32_core/pcpi_rs1$12$ , \picorv32_core/pcpi_rs2$12$ );  // ../src/picorv32.v(1232)
  and \picorv32_core/u117  (\picorv32_core/n443 [13], \picorv32_core/pcpi_rs1$13$ , \picorv32_core/pcpi_rs2$13$ );  // ../src/picorv32.v(1232)
  or \picorv32_core/u118  (\picorv32_core/n644 , \picorv32_core/decoded_rs2 [3], \picorv32_core/decoded_rs2 [4]);  // ../src/picorv32.v(1329)
  or \picorv32_core/u119  (\picorv32_core/n643 , \picorv32_core/decoded_rs2 [2], \picorv32_core/n644 );  // ../src/picorv32.v(1329)
  not \picorv32_core/u121  (\picorv32_core/n100 , \picorv32_core/n461 );  // ../src/picorv32.v(504)
  or \picorv32_core/u122  (\picorv32_core/n461 , \picorv32_core/n464 , \picorv32_core/n462 );  // ../src/picorv32.v(504)
  or \picorv32_core/u124  (\picorv32_core/n464 , \picorv32_core/n99 , \picorv32_core/n98 );  // ../src/picorv32.v(504)
  or \picorv32_core/u125  (\picorv32_core/n462 , \picorv32_core/n97 , \picorv32_core/n96 );  // ../src/picorv32.v(504)
  and \picorv32_core/u126  (\picorv32_core/n443 [14], \picorv32_core/pcpi_rs1$14$ , \picorv32_core/pcpi_rs2$14$ );  // ../src/picorv32.v(1232)
  or \picorv32_core/u127  (\picorv32_core/n101 , \picorv32_core/n99 , \picorv32_core/n462 );  // ../src/picorv32.v(504)
  and \picorv32_core/u128  (\picorv32_core/n443 [15], \picorv32_core/pcpi_rs1$15$ , \picorv32_core/pcpi_rs2$15$ );  // ../src/picorv32.v(1232)
  or \picorv32_core/u129  (\picorv32_core/n106 , \picorv32_core/n100 , \picorv32_core/n466 );  // ../src/picorv32.v(504)
  and \picorv32_core/u13  (\picorv32_core/mem_la_use_prefetched_high_word , \picorv32_core/n4 , \picorv32_core/clear_prefetched_high_word_neg );  // ../src/picorv32.v(336)
  and \picorv32_core/u130  (\picorv32_core/n443 [16], \picorv32_core/pcpi_rs1$16$ , \picorv32_core/pcpi_rs2$16$ );  // ../src/picorv32.v(1232)
  or \picorv32_core/u131  (\picorv32_core/n104 , \picorv32_core/n97 , \picorv32_core/n99 );  // ../src/picorv32.v(504)
  and \picorv32_core/u133  (\picorv32_core/n116 [3], mem_la_wstrb[3], mem_la_write);  // ../src/picorv32.v(540)
  or \picorv32_core/u134  (\picorv32_core/n675 , \picorv32_core/n668 , \picorv32_core/n686 );  // ../src/picorv32.v(1851)
  and \picorv32_core/u135  (\picorv32_core/n116 [2], mem_la_wstrb[2], mem_la_write);  // ../src/picorv32.v(540)
  or \picorv32_core/u136  (\picorv32_core/n680 , \picorv32_core/n666 , \picorv32_core/n662 );  // ../src/picorv32.v(1851)
  and \picorv32_core/u137  (\picorv32_core/n116 [1], mem_la_wstrb[1], mem_la_write);  // ../src/picorv32.v(540)
  or \picorv32_core/u138  (\picorv32_core/n670 , \picorv32_core/n684 , \picorv32_core/n680 );  // ../src/picorv32.v(1851)
  not \picorv32_core/u139  (\picorv32_core/n130 , \picorv32_core/n467 );  // ../src/picorv32.v(574)
  or \picorv32_core/u140  (\picorv32_core/n529 , \picorv32_core/is_slli_srli_srai , \picorv32_core/n448 );  // ../src/picorv32.v(1694)
  not \picorv32_core/u141  (\picorv32_core/instr_trap , \picorv32_core/n468 );  // ../src/picorv32.v(648)
  and \picorv32_core/u142  (\picorv32_core/n443 [17], \picorv32_core/pcpi_rs1$17$ , \picorv32_core/pcpi_rs2$17$ );  // ../src/picorv32.v(1232)
  or \picorv32_core/u143  (\picorv32_core/n468 , \picorv32_core/n492 , \picorv32_core/n469 );  // ../src/picorv32.v(648)
  or \picorv32_core/u144  (\picorv32_core/n458 , \picorv32_core/n645 , \picorv32_core/n643 );  // ../src/picorv32.v(1329)
  or \picorv32_core/u145  (\picorv32_core/n469 , \picorv32_core/n481 , \picorv32_core/n470 );  // ../src/picorv32.v(648)
  or \picorv32_core/u146  (\picorv32_core/n639 , \picorv32_core/decoded_rs1 [3], \picorv32_core/decoded_rs1 [4]);  // ../src/picorv32.v(1328)
  or \picorv32_core/u147  (\picorv32_core/n470 , \picorv32_core/n476 , \picorv32_core/n471 );  // ../src/picorv32.v(648)
  or \picorv32_core/u148  (\picorv32_core/n111 , \picorv32_core/n407 , trap);  // ../src/picorv32.v(530)
  and \picorv32_core/u15  (\picorv32_core/n7 , \picorv32_core/mem_la_use_prefetched_high_word , \picorv32_core/mem_do_rinst );  // ../src/picorv32.v(337)
  or \picorv32_core/u150  (\picorv32_core/n471 , \picorv32_core/n474 , \picorv32_core/n472 );  // ../src/picorv32.v(648)
  or \picorv32_core/u154  (\picorv32_core/n466 , \picorv32_core/n99 , \picorv32_core/n96 );  // ../src/picorv32.v(504)
  or \picorv32_core/u155  (\picorv32_core/n472 , \picorv32_core/instr_jal , \picorv32_core/n473 );  // ../src/picorv32.v(648)
  or \picorv32_core/u156  (\picorv32_core/n473 , \picorv32_core/instr_auipc , \picorv32_core/instr_lui );  // ../src/picorv32.v(648)
  or \picorv32_core/u157  (\picorv32_core/n474 , \picorv32_core/instr_bne , \picorv32_core/n475 );  // ../src/picorv32.v(648)
  or \picorv32_core/u158  (\picorv32_core/n475 , \picorv32_core/instr_beq , \picorv32_core/instr_jalr );  // ../src/picorv32.v(648)
  AL_MUX \picorv32_core/u159  (
    .i0(\picorv32_core/mem_valid ),
    .i1(\picorv32_core/mem_la_use_prefetched_high_word_neg ),
    .sel(\picorv32_core/n120 ),
    .o(\picorv32_core/n121 ));  // ../src/picorv32.v(552)
  or \picorv32_core/u16  (\picorv32_core/mem_xfer , \picorv32_core/mem_valid , \picorv32_core/n7 );  // ../src/picorv32.v(337)
  AL_MUX \picorv32_core/u161  (
    .i0(\picorv32_core/n121 ),
    .i1(1'b1),
    .sel(\picorv32_core/mem_do_wdata ),
    .o(\picorv32_core/n125 ));  // ../src/picorv32.v(557)
  not \picorv32_core/u164  (\picorv32_core/n598 , \picorv32_core/mem_do_rdata );  // ../src/picorv32.v(573)
  and \picorv32_core/u165  (\picorv32_core/n116 [0], mem_la_wstrb[0], mem_la_write);  // ../src/picorv32.v(540)
  or \picorv32_core/u166  (\picorv32_core/n131 , \picorv32_core/n130 , \picorv32_core/mem_la_secondword );  // ../src/picorv32.v(574)
  or \picorv32_core/u168  (\picorv32_core/n476 , \picorv32_core/n479 , \picorv32_core/n477 );  // ../src/picorv32.v(648)
  not \picorv32_core/u169  (\picorv32_core/n449 [2], \picorv32_core/latched_compr );  // ../src/picorv32.v(1270)
  and \picorv32_core/u170_sel_is_2  (\picorv32_core/u170_sel_is_2_o , \picorv32_core/mem_la_read_neg , \picorv32_core/n598 );
  AL_MUX \picorv32_core/u171  (
    .i0(\picorv32_core/mem_valid ),
    .i1(\picorv32_core/mem_la_read ),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n139 ));  // ../src/picorv32.v(583)
  and \picorv32_core/u173_sel_is_3  (\picorv32_core/u173_sel_is_3_o , \picorv32_core/mem_xfer , \picorv32_core/u170_sel_is_2_o );
  AL_MUX \picorv32_core/u174  (
    .i0(\picorv32_core/mem_valid ),
    .i1(1'b0),
    .sel(\picorv32_core/mem_xfer ),
    .o(\picorv32_core/n144 ));  // ../src/picorv32.v(591)
  and \picorv32_core/u179_sel_is_0  (\picorv32_core/u179_sel_is_0_o , \picorv32_core/clear_prefetched_high_word_neg , \picorv32_core/n111_neg );
  and \picorv32_core/u18  (\picorv32_core/n9 , \picorv32_core/mem_xfer , \picorv32_core/n8 );  // ../src/picorv32.v(340)
  and \picorv32_core/u180  (\picorv32_core/n467 , mem_rdata[0], mem_rdata[1]);  // ../src/picorv32.v(574)
  or \picorv32_core/u182  (\picorv32_core/n129 , \picorv32_core/instr_rdinstrh , \picorv32_core/instr_rdinstr );  // ../src/picorv32.v(651)
  or \picorv32_core/u184  (\picorv32_core/n607 , \picorv32_core/instr_add , \picorv32_core/instr_addi );  // ../src/picorv32.v(822)
  or \picorv32_core/u185  (\picorv32_core/n608 , \picorv32_core/instr_blt , \picorv32_core/instr_slti );  // ../src/picorv32.v(823)
  or \picorv32_core/u186  (\picorv32_core/n609 , \picorv32_core/instr_bltu , \picorv32_core/instr_sltiu );  // ../src/picorv32.v(824)
  or \picorv32_core/u187  (\picorv32_core/n610 , \picorv32_core/instr_lhu , \picorv32_core/instr_lbu );  // ../src/picorv32.v(825)
  and \picorv32_core/u188  (\picorv32_core/n170 , \picorv32_core/mem_do_rinst , \picorv32_core/mem_done );  // ../src/picorv32.v(828)
  or \picorv32_core/u189  (\picorv32_core/n613 , \picorv32_core/instr_sltu , \picorv32_core/instr_sltiu );  // ../src/picorv32.v(826)
  or \picorv32_core/u19  (\picorv32_core/n10 , \picorv32_core/mem_do_rinst , \picorv32_core/mem_do_rdata );  // ../src/picorv32.v(340)
  or \picorv32_core/u190  (\picorv32_core/n477 , \picorv32_core/instr_bltu , \picorv32_core/n478 );  // ../src/picorv32.v(648)
  or \picorv32_core/u191  (\picorv32_core/n478 , \picorv32_core/instr_bge , \picorv32_core/instr_blt );  // ../src/picorv32.v(648)
  or \picorv32_core/u192  (\picorv32_core/n479 , \picorv32_core/instr_lh , \picorv32_core/n480 );  // ../src/picorv32.v(648)
  or \picorv32_core/u193  (\picorv32_core/n619 , \picorv32_core/mem_rdata_latched [5], \picorv32_core/mem_rdata_latched [6]);  // ../src/picorv32.v(868)
  AL_MUX \picorv32_core/u194  (
    .i0(\picorv32_core/n178 ),
    .i1(\picorv32_core/n181 ),
    .sel(\picorv32_core/n96 ),
    .o(\picorv32_core/n183 ));  // ../src/picorv32.v(882)
  or \picorv32_core/u195  (\picorv32_core/n184 , \picorv32_core/n96 , \picorv32_core/n44 );  // ../src/picorv32.v(882)
  not \picorv32_core/u196  (\picorv32_core/n185 , \picorv32_core/n184 );  // ../src/picorv32.v(882)
  or \picorv32_core/u197  (\picorv32_core/n480 , \picorv32_core/instr_lb , \picorv32_core/instr_bgeu );  // ../src/picorv32.v(648)
  or \picorv32_core/u198  (\picorv32_core/n182 , \picorv32_core/n666 , \picorv32_core/n665 );  // ../src/picorv32.v(1851)
  or \picorv32_core/u199  (\picorv32_core/n481 , \picorv32_core/n487 , \picorv32_core/n482 );  // ../src/picorv32.v(648)
  or \picorv32_core/u20  (\picorv32_core/n11 , \picorv32_core/n10 , \picorv32_core/mem_do_wdata );  // ../src/picorv32.v(340)
  or \picorv32_core/u200  (\picorv32_core/n482 , \picorv32_core/n485 , \picorv32_core/n483 );  // ../src/picorv32.v(648)
  or \picorv32_core/u201  (\picorv32_core/n46 , \picorv32_core/n667 , \picorv32_core/n182 );  // ../src/picorv32.v(1851)
  or \picorv32_core/u202  (\picorv32_core/n188 , \picorv32_core/n96 , \picorv32_core/n97 );  // ../src/picorv32.v(882)
  or \picorv32_core/u203  (\picorv32_core/n483 , \picorv32_core/instr_lhu , \picorv32_core/n484 );  // ../src/picorv32.v(648)
  or \picorv32_core/u204  (\picorv32_core/n484 , \picorv32_core/instr_lbu , \picorv32_core/instr_lw );  // ../src/picorv32.v(648)
  or \picorv32_core/u205  (\picorv32_core/n48 , \picorv32_core/n663 , \picorv32_core/n662 );  // ../src/picorv32.v(1851)
  or \picorv32_core/u206  (\picorv32_core/n485 , \picorv32_core/instr_sw , \picorv32_core/n486 );  // ../src/picorv32.v(648)
  or \picorv32_core/u207  (\picorv32_core/n593 , \picorv32_core/n664 , \picorv32_core/n48 );  // ../src/picorv32.v(1851)
  AL_MUX \picorv32_core/u208  (
    .i0(\picorv32_core/n176 ),
    .i1(1'b1),
    .sel(\picorv32_core/n97 ),
    .o(\picorv32_core/n190 ));  // ../src/picorv32.v(882)
  AL_MUX \picorv32_core/u209  (
    .i0(\picorv32_core/n177 ),
    .i1(1'b1),
    .sel(\picorv32_core/n99 ),
    .o(\picorv32_core/n191 ));  // ../src/picorv32.v(882)
  and \picorv32_core/u21  (\picorv32_core/n12 , \picorv32_core/n9 , \picorv32_core/n11 );  // ../src/picorv32.v(340)
  or \picorv32_core/u210  (\picorv32_core/n486 , \picorv32_core/instr_sh , \picorv32_core/instr_sb );  // ../src/picorv32.v(648)
  AL_MUX \picorv32_core/u211  (
    .i0(\picorv32_core/n178 ),
    .i1(1'b1),
    .sel(\picorv32_core/n193 ),
    .o(\picorv32_core/n194 ));  // ../src/picorv32.v(909)
  not \picorv32_core/u213  (\picorv32_core/n197 , \picorv32_core/mem_rdata_latched [11]);  // ../src/picorv32.v(912)
  or \picorv32_core/u215  (\picorv32_core/n487 , \picorv32_core/n490 , \picorv32_core/n488 );  // ../src/picorv32.v(648)
  or \picorv32_core/u216  (\picorv32_core/n488 , \picorv32_core/instr_sltiu , \picorv32_core/n489 );  // ../src/picorv32.v(648)
  AL_MUX \picorv32_core/u217  (
    .i0(1'b1),
    .i1(\picorv32_core/n178 ),
    .sel(\picorv32_core/mux75_b0_sel_is_0_o ),
    .o(\picorv32_core/n201 ));
  or \picorv32_core/u218  (\picorv32_core/n489 , \picorv32_core/instr_slti , \picorv32_core/instr_addi );  // ../src/picorv32.v(648)
  or \picorv32_core/u219  (\picorv32_core/n490 , \picorv32_core/instr_andi , \picorv32_core/n491 );  // ../src/picorv32.v(648)
  or \picorv32_core/u22  (\picorv32_core/n8 , \picorv32_core/mem_state [0], \picorv32_core/mem_state [1]);  // ../src/picorv32.v(340)
  or \picorv32_core/u221  (\picorv32_core/n491 , \picorv32_core/instr_ori , \picorv32_core/instr_xori );  // ../src/picorv32.v(648)
  or \picorv32_core/u222  (\picorv32_core/n492 , \picorv32_core/n539 , \picorv32_core/n493 );  // ../src/picorv32.v(648)
  or \picorv32_core/u223  (\picorv32_core/n493 , \picorv32_core/n533 , \picorv32_core/n494 );  // ../src/picorv32.v(648)
  or \picorv32_core/u224  (\picorv32_core/n494 , \picorv32_core/n498 , \picorv32_core/n495 );  // ../src/picorv32.v(648)
  or \picorv32_core/u226  (\picorv32_core/n495 , \picorv32_core/instr_srai , \picorv32_core/n497 );  // ../src/picorv32.v(648)
  or \picorv32_core/u227  (\picorv32_core/n497 , \picorv32_core/instr_srli , \picorv32_core/instr_slli );  // ../src/picorv32.v(648)
  or \picorv32_core/u228  (\picorv32_core/n498 , \picorv32_core/instr_sll , \picorv32_core/n499 );  // ../src/picorv32.v(648)
  and \picorv32_core/u23  (\picorv32_core/n14 , \picorv32_core/n13 , \picorv32_core/mem_do_rinst );  // ../src/picorv32.v(340)
  or \picorv32_core/u230  (\picorv32_core/n499 , \picorv32_core/instr_sub , \picorv32_core/instr_add );  // ../src/picorv32.v(648)
  or \picorv32_core/u231  (\picorv32_core/n533 , \picorv32_core/n536 , \picorv32_core/n534 );  // ../src/picorv32.v(648)
  or \picorv32_core/u232  (\picorv32_core/n534 , \picorv32_core/instr_xor , \picorv32_core/n535 );  // ../src/picorv32.v(648)
  or \picorv32_core/u233  (\picorv32_core/n535 , \picorv32_core/instr_sltu , \picorv32_core/instr_slt );  // ../src/picorv32.v(648)
  or \picorv32_core/u234  (\picorv32_core/n536 , \picorv32_core/instr_or , \picorv32_core/n537 );  // ../src/picorv32.v(648)
  not \picorv32_core/u235_sel_is_0_o_inv  (\picorv32_core/u235_sel_is_0_o_neg , \picorv32_core/mux38_b0_sel_is_0_o );
  or \picorv32_core/u236  (\picorv32_core/n537 , \picorv32_core/instr_sra , \picorv32_core/instr_srl );  // ../src/picorv32.v(648)
  or \picorv32_core/u238  (\picorv32_core/n539 , \picorv32_core/n129 , \picorv32_core/n540 );  // ../src/picorv32.v(648)
  not \picorv32_core/u239_sel_is_0_o_inv  (\picorv32_core/u239_sel_is_0_o_neg , \picorv32_core/mux94_b0_sel_is_0_o );
  or \picorv32_core/u24  (\picorv32_core/n15 , \picorv32_core/n12 , \picorv32_core/n14 );  // ../src/picorv32.v(340)
  or \picorv32_core/u240  (\picorv32_core/n540 , \picorv32_core/instr_rdcycleh , \picorv32_core/n541 );  // ../src/picorv32.v(648)
  or \picorv32_core/u241  (\picorv32_core/n541 , \picorv32_core/instr_rdcycle , \picorv32_core/instr_and );  // ../src/picorv32.v(648)
  AL_MUX \picorv32_core/u245  (
    .i0(\picorv32_core/n178 ),
    .i1(1'b1),
    .sel(\picorv32_core/n96 ),
    .o(\picorv32_core/n228 ));  // ../src/picorv32.v(987)
  and \picorv32_core/u247_sel_is_1  (\picorv32_core/u247_sel_is_1_o , \picorv32_core/n98 , \picorv32_core/u235_sel_is_0_o_neg );
  AL_MUX \picorv32_core/u248  (
    .i0(\picorv32_core/n179 ),
    .i1(1'b1),
    .sel(\picorv32_core/u248_sel_is_1_o ),
    .o(\picorv32_core/n233 ));
  and \picorv32_core/u248_sel_is_1  (\picorv32_core/u248_sel_is_1_o , \picorv32_core/n98 , \picorv32_core/u239_sel_is_0_o_neg );
  and \picorv32_core/u25  (\picorv32_core/n16 , resetn, \picorv32_core/n15 );  // ../src/picorv32.v(340)
  AL_MUX \picorv32_core/u250  (
    .i0(\picorv32_core/n178 ),
    .i1(\picorv32_core/n234 ),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n249 ));  // ../src/picorv32.v(990)
  AL_MUX \picorv32_core/u251  (
    .i0(\picorv32_core/n176 ),
    .i1(\picorv32_core/n238 ),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n250 ));  // ../src/picorv32.v(990)
  AL_MUX \picorv32_core/u252  (
    .i0(\picorv32_core/n174 ),
    .i1(1'b1),
    .sel(\picorv32_core/u252_sel_is_3_o ),
    .o(\picorv32_core/n251 ));
  and \picorv32_core/u252_sel_is_3  (\picorv32_core/u252_sel_is_3_o , \picorv32_core/n180 , \picorv32_core/mux100_sel_is_6_o );
  AL_MUX \picorv32_core/u253  (
    .i0(\picorv32_core/n179 ),
    .i1(\picorv32_core/n240 ),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n252 ));  // ../src/picorv32.v(990)
  AL_MUX \picorv32_core/u254  (
    .i0(\picorv32_core/n177 ),
    .i1(\picorv32_core/n241 ),
    .sel(\picorv32_core/n180 ),
    .o(\picorv32_core/n253 ));  // ../src/picorv32.v(990)
  AL_MUX \picorv32_core/u255  (
    .i0(\picorv32_core/n175 ),
    .i1(1'b1),
    .sel(\picorv32_core/u255_sel_is_3_o ),
    .o(\picorv32_core/n254 ));
  and \picorv32_core/u255_sel_is_3  (\picorv32_core/u255_sel_is_3_o , \picorv32_core/n180 , \picorv32_core/mux103_sel_is_5_o );
  AL_MUX \picorv32_core/u256  (
    .i0(\picorv32_core/n173 ),
    .i1(1'b1),
    .sel(\picorv32_core/u256_sel_is_3_o ),
    .o(\picorv32_core/n255 ));
  and \picorv32_core/u256_sel_is_3  (\picorv32_core/u256_sel_is_3_o , \picorv32_core/n180 , \picorv32_core/mux104_sel_is_5_o );
  AL_MUX \picorv32_core/u257  (
    .i0(\picorv32_core/n171 ),
    .i1(1'b1),
    .sel(\picorv32_core/u257_sel_is_3_o ),
    .o(\picorv32_core/n256 ));
  and \picorv32_core/u257_sel_is_3  (\picorv32_core/u257_sel_is_3_o , \picorv32_core/n180 , \picorv32_core/mux105_sel_is_5_o );
  and \picorv32_core/u27  (\picorv32_core/n13 , \picorv32_core/mem_state [0], \picorv32_core/mem_state [1]);  // ../src/picorv32.v(340)
  not \picorv32_core/u270  (\picorv32_core/n273 , \picorv32_core/decoder_pseudo_trigger );  // ../src/picorv32.v(993)
  and \picorv32_core/u271  (\picorv32_core/n274 , \picorv32_core/decoder_trigger , \picorv32_core/n273 );  // ../src/picorv32.v(993)
  and \picorv32_core/u272  (\picorv32_core/n276 , \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu , \picorv32_core/n275 );  // ../src/picorv32.v(996)
  and \picorv32_core/u273  (\picorv32_core/n278 , \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu , \picorv32_core/n277 );  // ../src/picorv32.v(997)
  and \picorv32_core/u274  (\picorv32_core/n280 , \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu , \picorv32_core/n279 );  // ../src/picorv32.v(998)
  and \picorv32_core/u275  (\picorv32_core/n282 , \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu , \picorv32_core/n281 );  // ../src/picorv32.v(999)
  and \picorv32_core/u276  (\picorv32_core/n284 , \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu , \picorv32_core/n283 );  // ../src/picorv32.v(1000)
  and \picorv32_core/u277  (\picorv32_core/n286 , \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu , \picorv32_core/n285 );  // ../src/picorv32.v(1001)
  or \picorv32_core/u278  (\picorv32_core/is_rdcycle_rdcycleh_rdinstr_rdinstrh , \picorv32_core/n129 , \picorv32_core/n573 );  // ../src/picorv32.v(651)
  and \picorv32_core/u279  (\picorv32_core/n287 , \picorv32_core/is_lb_lh_lw_lbu_lhu , \picorv32_core/n275 );  // ../src/picorv32.v(1003)
  and \picorv32_core/u28  (\picorv32_core/n19 , \picorv32_core/n18 , \picorv32_core/mem_xfer );  // ../src/picorv32.v(341)
  or \picorv32_core/u280  (\picorv32_core/n573 , \picorv32_core/instr_rdcycleh , \picorv32_core/instr_rdcycle );  // ../src/picorv32.v(651)
  and \picorv32_core/u281  (\picorv32_core/n288 , \picorv32_core/is_lb_lh_lw_lbu_lhu , \picorv32_core/n277 );  // ../src/picorv32.v(1004)
  and \picorv32_core/u282  (\picorv32_core/n290 , \picorv32_core/is_lb_lh_lw_lbu_lhu , \picorv32_core/n289 );  // ../src/picorv32.v(1005)
  and \picorv32_core/u284  (\picorv32_core/n291 , \picorv32_core/is_lb_lh_lw_lbu_lhu , \picorv32_core/n279 );  // ../src/picorv32.v(1006)
  or \picorv32_core/u285  (\picorv32_core/n165 , \picorv32_core/n606 , \picorv32_core/n603 );  // ../src/picorv32.v(822)
  and \picorv32_core/u286  (\picorv32_core/n292 , \picorv32_core/is_lb_lh_lw_lbu_lhu , \picorv32_core/n281 );  // ../src/picorv32.v(1007)
  or \picorv32_core/u287  (\picorv32_core/n603 , \picorv32_core/n605 , \picorv32_core/n473 );  // ../src/picorv32.v(822)
  and \picorv32_core/u288  (\picorv32_core/n293 , \picorv32_core/is_sb_sh_sw , \picorv32_core/n275 );  // ../src/picorv32.v(1009)
  or \picorv32_core/u29  (\picorv32_core/n20 , \picorv32_core/mem_la_firstword_neg , \picorv32_core/n19 );  // ../src/picorv32.v(341)
  and \picorv32_core/u290  (\picorv32_core/n294 , \picorv32_core/is_sb_sh_sw , \picorv32_core/n277 );  // ../src/picorv32.v(1010)
  or \picorv32_core/u291  (\picorv32_core/n605 , \picorv32_core/instr_jalr , \picorv32_core/instr_jal );  // ../src/picorv32.v(822)
  and \picorv32_core/u292  (\picorv32_core/n295 , \picorv32_core/is_sb_sh_sw , \picorv32_core/n289 );  // ../src/picorv32.v(1011)
  or \picorv32_core/u293  (\picorv32_core/n606 , \picorv32_core/instr_sub , \picorv32_core/n607 );  // ../src/picorv32.v(822)
  and \picorv32_core/u294  (\picorv32_core/n296 , \picorv32_core/is_alu_reg_imm , \picorv32_core/n275 );  // ../src/picorv32.v(1013)
  or \picorv32_core/u295  (\picorv32_core/n166 , \picorv32_core/instr_slt , \picorv32_core/n608 );  // ../src/picorv32.v(823)
  and \picorv32_core/u296  (\picorv32_core/n297 , \picorv32_core/is_alu_reg_imm , \picorv32_core/n289 );  // ../src/picorv32.v(1014)
  and \picorv32_core/u297  (\picorv32_core/n299 , \picorv32_core/is_alu_reg_imm , \picorv32_core/n298 );  // ../src/picorv32.v(1015)
  or \picorv32_core/u298  (\picorv32_core/n167 , \picorv32_core/instr_sltu , \picorv32_core/n609 );  // ../src/picorv32.v(824)
  and \picorv32_core/u299  (\picorv32_core/n300 , \picorv32_core/is_alu_reg_imm , \picorv32_core/n279 );  // ../src/picorv32.v(1016)
  and \picorv32_core/u30  (\picorv32_core/mem_done , \picorv32_core/n16 , \picorv32_core/n20 );  // ../src/picorv32.v(341)
  or \picorv32_core/u300  (\picorv32_core/n168 , \picorv32_core/instr_lw , \picorv32_core/n610 );  // ../src/picorv32.v(825)
  and \picorv32_core/u301  (\picorv32_core/n301 , \picorv32_core/is_alu_reg_imm , \picorv32_core/n283 );  // ../src/picorv32.v(1017)
  or \picorv32_core/u302  (\picorv32_core/n169 , \picorv32_core/n613 , \picorv32_core/n611 );  // ../src/picorv32.v(826)
  and \picorv32_core/u303  (\picorv32_core/n302 , \picorv32_core/is_alu_reg_imm , \picorv32_core/n285 );  // ../src/picorv32.v(1018)
  or \picorv32_core/u304  (\picorv32_core/n611 , \picorv32_core/instr_slt , \picorv32_core/n612 );  // ../src/picorv32.v(826)
  and \picorv32_core/u305  (\picorv32_core/n303 , \picorv32_core/is_alu_reg_imm , \picorv32_core/n277 );  // ../src/picorv32.v(1020)
  and \picorv32_core/u306  (\picorv32_core/n305 , \picorv32_core/n303 , \picorv32_core/n304 );  // ../src/picorv32.v(1020)
  or \picorv32_core/u307  (\picorv32_core/n612 , \picorv32_core/instr_slti , \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );  // ../src/picorv32.v(826)
  and \picorv32_core/u308  (\picorv32_core/n306 , \picorv32_core/is_alu_reg_imm , \picorv32_core/n281 );  // ../src/picorv32.v(1021)
  or \picorv32_core/u309  (\picorv32_core/n181 , \picorv32_core/n617 , \picorv32_core/n614 );  // ../src/picorv32.v(868)
  and \picorv32_core/u31  (\picorv32_core/n351 , \picorv32_core/mem_rdata_latched [0], \picorv32_core/mem_rdata_latched [1]);  // ../src/picorv32.v(341)
  and \picorv32_core/u310  (\picorv32_core/n307 , \picorv32_core/n306 , \picorv32_core/n304 );  // ../src/picorv32.v(1021)
  or \picorv32_core/u311  (\picorv32_core/n614 , \picorv32_core/n616 , \picorv32_core/n615 );  // ../src/picorv32.v(868)
  or \picorv32_core/u312  (\picorv32_core/n615 , \picorv32_core/mem_rdata_latched [11], \picorv32_core/mem_rdata_latched [12]);  // ../src/picorv32.v(868)
  and \picorv32_core/u313  (\picorv32_core/n309 , \picorv32_core/n306 , \picorv32_core/n308 );  // ../src/picorv32.v(1022)
  or \picorv32_core/u314  (\picorv32_core/n616 , \picorv32_core/mem_rdata_latched [9], \picorv32_core/mem_rdata_latched [10]);  // ../src/picorv32.v(868)
  and \picorv32_core/u315  (\picorv32_core/n310 , \picorv32_core/is_alu_reg_reg , \picorv32_core/n275 );  // ../src/picorv32.v(1024)
  or \picorv32_core/u316  (\picorv32_core/n617 , \picorv32_core/n619 , \picorv32_core/n618 );  // ../src/picorv32.v(868)
  and \picorv32_core/u317  (\picorv32_core/n311 , \picorv32_core/n310 , \picorv32_core/n304 );  // ../src/picorv32.v(1024)
  or \picorv32_core/u318  (\picorv32_core/n618 , \picorv32_core/mem_rdata_latched [7], \picorv32_core/mem_rdata_latched [8]);  // ../src/picorv32.v(868)
  not \picorv32_core/u319  (\picorv32_core/n44 , \picorv32_core/n101 );  // ../src/picorv32.v(882)
  and \picorv32_core/u32  (\picorv32_core/n22 , resetn, \picorv32_core/n21 );  // ../src/picorv32.v(343)
  and \picorv32_core/u321  (\picorv32_core/n312 , \picorv32_core/n310 , \picorv32_core/n308 );  // ../src/picorv32.v(1025)
  or \picorv32_core/u322  (\picorv32_core/n346 , \picorv32_core/n345 , \picorv32_core/n622 );  // ../src/picorv32.v(1054)
  and \picorv32_core/u323  (\picorv32_core/n313 , \picorv32_core/is_alu_reg_reg , \picorv32_core/n277 );  // ../src/picorv32.v(1026)
  or \picorv32_core/u324  (\picorv32_core/n348 , \picorv32_core/n625 , \picorv32_core/n623 );  // ../src/picorv32.v(1063)
  and \picorv32_core/u325  (\picorv32_core/n314 , \picorv32_core/n313 , \picorv32_core/n304 );  // ../src/picorv32.v(1026)
  or \picorv32_core/u326  (\picorv32_core/n623 , \picorv32_core/n298 , \picorv32_core/n624 );  // ../src/picorv32.v(1063)
  and \picorv32_core/u327  (\picorv32_core/n315 , \picorv32_core/is_alu_reg_reg , \picorv32_core/n289 );  // ../src/picorv32.v(1027)
  or \picorv32_core/u328  (\picorv32_core/n624 , \picorv32_core/n289 , \picorv32_core/n275 );  // ../src/picorv32.v(1063)
  and \picorv32_core/u329  (\picorv32_core/n316 , \picorv32_core/n315 , \picorv32_core/n304 );  // ../src/picorv32.v(1027)
  and \picorv32_core/u33  (mem_la_write, \picorv32_core/n22 , \picorv32_core/mem_do_wdata );  // ../src/picorv32.v(343)
  or \picorv32_core/u330  (\picorv32_core/n625 , \picorv32_core/n285 , \picorv32_core/n626 );  // ../src/picorv32.v(1063)
  and \picorv32_core/u331  (\picorv32_core/n317 , \picorv32_core/is_alu_reg_reg , \picorv32_core/n298 );  // ../src/picorv32.v(1028)
  or \picorv32_core/u332  (\picorv32_core/n356 , \picorv32_core/is_alu_reg_imm , \picorv32_core/n627 );  // ../src/picorv32.v(1080)
  and \picorv32_core/u333  (\picorv32_core/n318 , \picorv32_core/n317 , \picorv32_core/n304 );  // ../src/picorv32.v(1028)
  and \picorv32_core/u335  (\picorv32_core/n319 , \picorv32_core/is_alu_reg_reg , \picorv32_core/n279 );  // ../src/picorv32.v(1029)
  and \picorv32_core/u337  (\picorv32_core/n320 , \picorv32_core/n319 , \picorv32_core/n304 );  // ../src/picorv32.v(1029)
  and \picorv32_core/u339  (\picorv32_core/n321 , \picorv32_core/is_alu_reg_reg , \picorv32_core/n281 );  // ../src/picorv32.v(1030)
  and \picorv32_core/u341  (\picorv32_core/n322 , \picorv32_core/n321 , \picorv32_core/n304 );  // ../src/picorv32.v(1030)
  xor \picorv32_core/u342  (\picorv32_core/n439 [31], \picorv32_core/pcpi_rs1$31$ , \picorv32_core/pcpi_rs2$31$ );  // ../src/picorv32.v(1228)
  xor \picorv32_core/u343  (\picorv32_core/n439 [30], \picorv32_core/pcpi_rs1$30$ , \picorv32_core/pcpi_rs2$30$ );  // ../src/picorv32.v(1228)
  xor \picorv32_core/u344  (\picorv32_core/n439 [29], \picorv32_core/pcpi_rs1$29$ , \picorv32_core/pcpi_rs2$29$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u345  (\picorv32_core/n323 , \picorv32_core/n321 , \picorv32_core/n308 );  // ../src/picorv32.v(1031)
  xor \picorv32_core/u346  (\picorv32_core/n439 [28], \picorv32_core/pcpi_rs1$28$ , \picorv32_core/pcpi_rs2$28$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u347  (\picorv32_core/n324 , \picorv32_core/is_alu_reg_reg , \picorv32_core/n283 );  // ../src/picorv32.v(1032)
  xor \picorv32_core/u348  (\picorv32_core/n439 [27], \picorv32_core/pcpi_rs1$27$ , \picorv32_core/pcpi_rs2$27$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u349  (\picorv32_core/n325 , \picorv32_core/n324 , \picorv32_core/n304 );  // ../src/picorv32.v(1032)
  xor \picorv32_core/u350  (\picorv32_core/n439 [26], \picorv32_core/pcpi_rs1$26$ , \picorv32_core/pcpi_rs2$26$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u351  (\picorv32_core/n326 , \picorv32_core/is_alu_reg_reg , \picorv32_core/n285 );  // ../src/picorv32.v(1033)
  xor \picorv32_core/u352  (\picorv32_core/n439 [25], \picorv32_core/pcpi_rs1$25$ , \picorv32_core/pcpi_rs2$25$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u353  (\picorv32_core/n327 , \picorv32_core/n326 , \picorv32_core/n304 );  // ../src/picorv32.v(1033)
  and \picorv32_core/u354  (\picorv32_core/n330 , \picorv32_core/n328 , \picorv32_core/n329 );  // ../src/picorv32.v(1035)
  xor \picorv32_core/u355  (\picorv32_core/n439 [24], \picorv32_core/pcpi_rs1$24$ , \picorv32_core/pcpi_rs2$24$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u356  (\picorv32_core/n332 , \picorv32_core/n328 , \picorv32_core/n331 );  // ../src/picorv32.v(1036)
  or \picorv32_core/u357  (\picorv32_core/n333 , \picorv32_core/n330 , \picorv32_core/n332 );  // ../src/picorv32.v(1036)
  xor \picorv32_core/u358  (\picorv32_core/n439 [23], \picorv32_core/pcpi_rs1$23$ , \picorv32_core/pcpi_rs2$23$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u359  (\picorv32_core/n335 , \picorv32_core/n328 , \picorv32_core/n334 );  // ../src/picorv32.v(1037)
  and \picorv32_core/u36  (\picorv32_core/n24 , \picorv32_core/mem_la_use_prefetched_high_word_neg , \picorv32_core/n21 );  // ../src/picorv32.v(344)
  xor \picorv32_core/u360  (\picorv32_core/n439 [22], \picorv32_core/pcpi_rs1$22$ , \picorv32_core/pcpi_rs2$22$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u361  (\picorv32_core/n337 , \picorv32_core/n328 , \picorv32_core/n336 );  // ../src/picorv32.v(1038)
  or \picorv32_core/u362  (\picorv32_core/n338 , \picorv32_core/n335 , \picorv32_core/n337 );  // ../src/picorv32.v(1038)
  xor \picorv32_core/u363  (\picorv32_core/n439 [21], \picorv32_core/pcpi_rs1$21$ , \picorv32_core/pcpi_rs2$21$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u364  (\picorv32_core/n340 , \picorv32_core/n328 , \picorv32_core/n339 );  // ../src/picorv32.v(1039)
  xor \picorv32_core/u365  (\picorv32_core/n439 [20], \picorv32_core/pcpi_rs1$20$ , \picorv32_core/pcpi_rs2$20$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u366  (\picorv32_core/n342 , \picorv32_core/n328 , \picorv32_core/n341 );  // ../src/picorv32.v(1040)
  xor \picorv32_core/u367  (\picorv32_core/n439 [19], \picorv32_core/pcpi_rs1$19$ , \picorv32_core/pcpi_rs2$19$ );  // ../src/picorv32.v(1228)
  xor \picorv32_core/u368  (\picorv32_core/n439 [18], \picorv32_core/pcpi_rs1$18$ , \picorv32_core/pcpi_rs2$18$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u369  (\picorv32_core/n343 , \picorv32_core/n277 , \picorv32_core/n304 );  // ../src/picorv32.v(1051)
  xor \picorv32_core/u370  (\picorv32_core/n439 [17], \picorv32_core/pcpi_rs1$17$ , \picorv32_core/pcpi_rs2$17$ );  // ../src/picorv32.v(1228)
  xor \picorv32_core/u371  (\picorv32_core/n439 [16], \picorv32_core/pcpi_rs1$16$ , \picorv32_core/pcpi_rs2$16$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u372  (\picorv32_core/n344 , \picorv32_core/n281 , \picorv32_core/n304 );  // ../src/picorv32.v(1052)
  xor \picorv32_core/u373  (\picorv32_core/n439 [15], \picorv32_core/pcpi_rs1$15$ , \picorv32_core/pcpi_rs2$15$ );  // ../src/picorv32.v(1228)
  xor \picorv32_core/u374  (\picorv32_core/n439 [14], \picorv32_core/pcpi_rs1$14$ , \picorv32_core/pcpi_rs2$14$ );  // ../src/picorv32.v(1228)
  and \picorv32_core/u375  (\picorv32_core/n345 , \picorv32_core/n281 , \picorv32_core/n308 );  // ../src/picorv32.v(1053)
  and \picorv32_core/u377  (\picorv32_core/n347 , \picorv32_core/is_alu_reg_imm , \picorv32_core/n346 );  // ../src/picorv32.v(1054)
  xor \picorv32_core/u378  (\picorv32_core/n439 [13], \picorv32_core/pcpi_rs1$13$ , \picorv32_core/pcpi_rs2$13$ );  // ../src/picorv32.v(1228)
  xor \picorv32_core/u379  (\picorv32_core/n439 [12], \picorv32_core/pcpi_rs1$12$ , \picorv32_core/pcpi_rs2$12$ );  // ../src/picorv32.v(1228)
  or \picorv32_core/u38  (\picorv32_core/n120 , \picorv32_core/n0 , \picorv32_core/mem_do_rdata );  // ../src/picorv32.v(344)
  xor \picorv32_core/u380  (\picorv32_core/n439 [11], \picorv32_core/pcpi_rs1$11$ , \picorv32_core/pcpi_rs2$11$ );  // ../src/picorv32.v(1228)
  xor \picorv32_core/u381  (\picorv32_core/n439 [10], \picorv32_core/pcpi_rs1$10$ , \picorv32_core/pcpi_rs2$10$ );  // ../src/picorv32.v(1228)
  xor \picorv32_core/u382  (\picorv32_core/n439 [9], \picorv32_core/pcpi_rs1$9$ , \picorv32_core/pcpi_rs2$9$ );  // ../src/picorv32.v(1228)
  xor \picorv32_core/u383  (\picorv32_core/n439 [8], \picorv32_core/pcpi_rs1$8$ , \picorv32_core/pcpi_rs2$8$ );  // ../src/picorv32.v(1228)
  or \picorv32_core/u384  (\picorv32_core/n622 , \picorv32_core/n344 , \picorv32_core/n343 );  // ../src/picorv32.v(1054)
  and \picorv32_core/u385  (\picorv32_core/n349 , \picorv32_core/is_alu_reg_imm , \picorv32_core/n348 );  // ../src/picorv32.v(1063)
  or \picorv32_core/u386  (\picorv32_core/n350 , \picorv32_core/instr_jalr , \picorv32_core/n349 );  // ../src/picorv32.v(1063)
  xor \picorv32_core/u387  (\picorv32_core/n439 [7], \picorv32_core/pcpi_rs1$7$ , mem_la_wdata[7]);  // ../src/picorv32.v(1228)
  xor \picorv32_core/u388  (\picorv32_core/n439 [6], \picorv32_core/pcpi_rs1$6$ , mem_la_wdata[6]);  // ../src/picorv32.v(1228)
  xor \picorv32_core/u389  (\picorv32_core/n439 [5], \picorv32_core/pcpi_rs1$5$ , mem_la_wdata[5]);  // ../src/picorv32.v(1228)
  and \picorv32_core/u39  (\picorv32_core/n25 , \picorv32_core/n24 , \picorv32_core/n120 );  // ../src/picorv32.v(344)
  xor \picorv32_core/u390  (\picorv32_core/n439 [4], \picorv32_core/pcpi_rs1$4$ , mem_la_wdata[4]);  // ../src/picorv32.v(1228)
  xor \picorv32_core/u391  (\picorv32_core/n439 [3], \picorv32_core/pcpi_rs1$3$ , mem_la_wdata[3]);  // ../src/picorv32.v(1228)
  xor \picorv32_core/u392  (\picorv32_core/n439 [2], \picorv32_core/pcpi_rs1$2$ , mem_la_wdata[2]);  // ../src/picorv32.v(1228)
  xor \picorv32_core/u393  (\picorv32_core/n439 [1], \picorv32_core/pcpi_rs1$1$ , mem_la_wdata[1]);  // ../src/picorv32.v(1228)
  or \picorv32_core/u394  (\picorv32_core/n441 [31], \picorv32_core/pcpi_rs1$31$ , \picorv32_core/pcpi_rs2$31$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u395  (\picorv32_core/n441 [30], \picorv32_core/pcpi_rs1$30$ , \picorv32_core/pcpi_rs2$30$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u396  (\picorv32_core/n441 [29], \picorv32_core/pcpi_rs1$29$ , \picorv32_core/pcpi_rs2$29$ );  // ../src/picorv32.v(1230)
  and \picorv32_core/u397  (\picorv32_core/n354 , \picorv32_core/is_alu_reg_reg , \picorv32_core/n346 );  // ../src/picorv32.v(1069)
  or \picorv32_core/u398  (\picorv32_core/n626 , \picorv32_core/n283 , \picorv32_core/n279 );  // ../src/picorv32.v(1063)
  or \picorv32_core/u4  (\picorv32_core/n0 , \picorv32_core/mem_do_prefetch , \picorv32_core/mem_do_rinst );  // ../src/picorv32.v(326)
  or \picorv32_core/u400  (\picorv32_core/n627 , \picorv32_core/is_lb_lh_lw_lbu_lhu , \picorv32_core/instr_jalr );  // ../src/picorv32.v(1080)
  and \picorv32_core/u44  (\picorv32_core/n26 , \picorv32_core/mem_la_firstword_xfer , \picorv32_core/mem_la_secondword_neg );  // ../src/picorv32.v(345)
  or \picorv32_core/u447  (\picorv32_core/n441 [28], \picorv32_core/pcpi_rs1$28$ , \picorv32_core/pcpi_rs2$28$ );  // ../src/picorv32.v(1230)
  and \picorv32_core/u449_sel_is_0  (\picorv32_core/u449_sel_is_0_o , resetn, \picorv32_core/n274_neg );
  and \picorv32_core/u46  (\picorv32_core/n28 , \picorv32_core/n26 , \picorv32_core/n351 );  // ../src/picorv32.v(345)
  or \picorv32_core/u47  (\picorv32_core/n29 , \picorv32_core/n25 , \picorv32_core/n28 );  // ../src/picorv32.v(345)
  and \picorv32_core/u472  (\picorv32_core/n432 , \picorv32_core/latched_store , \picorv32_core/latched_branch );  // ../src/picorv32.v(1166)
  not \picorv32_core/u474  (\picorv32_core/n436 , \picorv32_core/alu_lts );  // ../src/picorv32.v(1211)
  not \picorv32_core/u475  (\picorv32_core/n437 , \picorv32_core/alu_ltu );  // ../src/picorv32.v(1213)
  or \picorv32_core/u476  (\picorv32_core/n438 , \picorv32_core/instr_xori , \picorv32_core/instr_xor );  // ../src/picorv32.v(1227)
  or \picorv32_core/u478  (\picorv32_core/n440 , \picorv32_core/instr_ori , \picorv32_core/instr_or );  // ../src/picorv32.v(1229)
  xor \picorv32_core/u479  (\picorv32_core/n439 [0], \picorv32_core/pcpi_rs1$0$ , mem_la_wdata[0]);  // ../src/picorv32.v(1228)
  and \picorv32_core/u48  (\picorv32_core/mem_la_read , resetn, \picorv32_core/n29 );  // ../src/picorv32.v(345)
  or \picorv32_core/u480  (\picorv32_core/n442 , \picorv32_core/instr_andi , \picorv32_core/instr_and );  // ../src/picorv32.v(1231)
  or \picorv32_core/u481  (\picorv32_core/n441 [0], \picorv32_core/pcpi_rs1$0$ , mem_la_wdata[0]);  // ../src/picorv32.v(1230)
  AL_MUX \picorv32_core/u483  (
    .i0(1'b0),
    .i1(\picorv32_core/clear_prefetched_high_word_q ),
    .sel(\picorv32_core/prefetched_high_word ),
    .o(\picorv32_core/n444 ));  // ../src/picorv32.v(1246)
  and \picorv32_core/u484  (\picorv32_core/n443 [0], \picorv32_core/pcpi_rs1$0$ , mem_la_wdata[0]);  // ../src/picorv32.v(1232)
  or \picorv32_core/u486  (\picorv32_core/n441 [27], \picorv32_core/pcpi_rs1$27$ , \picorv32_core/pcpi_rs2$27$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u487  (\picorv32_core/n447 , \picorv32_core/latched_branch , \picorv32_core/n407 );  // ../src/picorv32.v(1247)
  AL_MUX \picorv32_core/u488  (
    .i0(\picorv32_core/n444 ),
    .i1(1'b1),
    .sel(\picorv32_core/n447 ),
    .o(\picorv32_core/clear_prefetched_high_word ));  // ../src/picorv32.v(1248)
  not \picorv32_core/u489  (\picorv32_core/n501 [2], \picorv32_core/compressed_instr );  // ../src/picorv32.v(1498)
  not \picorv32_core/u490  (\picorv32_core/n451 , \picorv32_core/latched_branch );  // ../src/picorv32.v(1273)
  and \picorv32_core/u491  (\picorv32_core/n452 , \picorv32_core/latched_store , \picorv32_core/n451 );  // ../src/picorv32.v(1273)
  AL_MUX \picorv32_core/u493  (
    .i0(1'b0),
    .i1(\picorv32_core/n632 ),
    .sel(\picorv32_core/n663 ),
    .o(\picorv32_core/cpuregs_write ));  // ../src/picorv32.v(1286)
  and \picorv32_core/u494  (\picorv32_core/n456 , \picorv32_core/cpuregs_write , resetn);  // ../src/picorv32.v(1313)
  or \picorv32_core/u495  (\picorv32_core/n441 [26], \picorv32_core/pcpi_rs1$26$ , \picorv32_core/pcpi_rs2$26$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u496  (\picorv32_core/n632 , \picorv32_core/n452 , \picorv32_core/latched_branch );  // ../src/picorv32.v(1285)
  or \picorv32_core/u497  (\picorv32_core/n640 , \picorv32_core/decoded_rs1 [0], \picorv32_core/decoded_rs1 [1]);  // ../src/picorv32.v(1328)
  or \picorv32_core/u498  (\picorv32_core/n441 [25], \picorv32_core/pcpi_rs1$25$ , \picorv32_core/pcpi_rs2$25$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u499  (\picorv32_core/n441 [24], \picorv32_core/pcpi_rs1$24$ , \picorv32_core/pcpi_rs2$24$ );  // ../src/picorv32.v(1230)
  and \picorv32_core/u5  (\picorv32_core/n1 , \picorv32_core/n0 , \picorv32_core/next_pc [1]);  // ../src/picorv32.v(326)
  not \picorv32_core/u50  (\picorv32_core/n407 , resetn);  // ../src/picorv32.v(355)
  not \picorv32_core/u500  (\picorv32_core/n463 , \picorv32_core/decoder_trigger );  // ../src/picorv32.v(1430)
  or \picorv32_core/u503  (\picorv32_core/n441 [23], \picorv32_core/pcpi_rs1$23$ , \picorv32_core/pcpi_rs2$23$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u504  (\picorv32_core/n441 [22], \picorv32_core/pcpi_rs1$22$ , \picorv32_core/pcpi_rs2$22$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u505  (\picorv32_core/n441 [21], \picorv32_core/pcpi_rs1$21$ , \picorv32_core/pcpi_rs2$21$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u506  (\picorv32_core/n441 [20], \picorv32_core/pcpi_rs1$20$ , \picorv32_core/pcpi_rs2$20$ );  // ../src/picorv32.v(1230)
  not \picorv32_core/u508  (\picorv32_core/n505 , \picorv32_core/instr_jalr );  // ../src/picorv32.v(1511)
  AL_MUX \picorv32_core/u512  (
    .i0(\picorv32_core/n463 ),
    .i1(\picorv32_core/instr_jal ),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n513 ));  // ../src/picorv32.v(1514)
  AL_MUX \picorv32_core/u513  (
    .i0(1'b0),
    .i1(\picorv32_core/instr_jal ),
    .sel(\picorv32_core/decoder_trigger ),
    .o(\picorv32_core/n514 ));  // ../src/picorv32.v(1514)
  and \picorv32_core/u515  (\picorv32_core/n519 , \picorv32_core/is_lb_lh_lw_lbu_lhu , \picorv32_core/n468 );  // ../src/picorv32.v(1634)
  or \picorv32_core/u516  (\picorv32_core/n645 , \picorv32_core/decoded_rs2 [0], \picorv32_core/decoded_rs2 [1]);  // ../src/picorv32.v(1329)
  or \picorv32_core/u517  (\picorv32_core/n646 , \picorv32_core/is_sll_srl_sra , \picorv32_core/is_sb_sh_sw );  // ../src/picorv32.v(1690)
  AL_MUX \picorv32_core/u518  (
    .i0(\picorv32_core/latched_store ),
    .i1(1'b1),
    .sel(\picorv32_core/is_rdcycle_rdcycleh_rdinstr_rdinstrh ),
    .o(\picorv32_core/n526 ));  // ../src/picorv32.v(1694)
  or \picorv32_core/u519  (\picorv32_core/n651 , \picorv32_core/is_slli_srli_srai , \picorv32_core/n519 );  // ../src/picorv32.v(1694)
  not \picorv32_core/u52  (\picorv32_core/n18 , \picorv32_core/n351 );  // ../src/picorv32.v(341)
  or \picorv32_core/u520  (\picorv32_core/n530 , \picorv32_core/is_lui_auipc_jal , \picorv32_core/is_jalr_addi_slti_sltiu_xori_ori_andi );  // ../src/picorv32.v(1694)
  or \picorv32_core/u521  (\picorv32_core/n441 [19], \picorv32_core/pcpi_rs1$19$ , \picorv32_core/pcpi_rs2$19$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u522  (\picorv32_core/n441 [18], \picorv32_core/pcpi_rs1$18$ , \picorv32_core/pcpi_rs2$18$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u523  (\picorv32_core/n441 [17], \picorv32_core/pcpi_rs1$17$ , \picorv32_core/pcpi_rs2$17$ );  // ../src/picorv32.v(1230)
  AL_MUX \picorv32_core/u525  (
    .i0(1'b1),
    .i1(\picorv32_core/alu_out_0 ),
    .sel(\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ),
    .o(\picorv32_core/n547 ));  // ../src/picorv32.v(1764)
  AL_MUX \picorv32_core/u526  (
    .i0(\picorv32_core/instr_jalr ),
    .i1(\picorv32_core/alu_out_0 ),
    .sel(\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ),
    .o(\picorv32_core/n548 ));  // ../src/picorv32.v(1764)
  AL_MUX \picorv32_core/u527  (
    .i0(\picorv32_core/n170 ),
    .i1(1'b0),
    .sel(\picorv32_core/u527_sel_is_3_o ),
    .o(\picorv32_core/n550 ));
  and \picorv32_core/u527_sel_is_3  (\picorv32_core/u527_sel_is_3_o , \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu , \picorv32_core/alu_out_0 );
  AL_MUX \picorv32_core/u529  (
    .i0(1'b1),
    .i1(\picorv32_core/latched_stalu ),
    .sel(\picorv32_core/is_beq_bne_blt_bge_bltu_bgeu ),
    .o(\picorv32_core/n552 ));  // ../src/picorv32.v(1764)
  or \picorv32_core/u530  (\picorv32_core/n555 , \picorv32_core/instr_slli , \picorv32_core/instr_sll );  // ../src/picorv32.v(1776)
  or \picorv32_core/u532  (\picorv32_core/n557 , \picorv32_core/instr_srai , \picorv32_core/instr_sra );  // ../src/picorv32.v(1778)
  and \picorv32_core/u533  (\picorv32_core/n443 [24], \picorv32_core/pcpi_rs1$24$ , \picorv32_core/pcpi_rs2$24$ );  // ../src/picorv32.v(1232)
  or \picorv32_core/u534  (\picorv32_core/n441 [16], \picorv32_core/pcpi_rs1$16$ , \picorv32_core/pcpi_rs2$16$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u535  (\picorv32_core/n441 [15], \picorv32_core/pcpi_rs1$15$ , \picorv32_core/pcpi_rs2$15$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u536  (\picorv32_core/n441 [14], \picorv32_core/pcpi_rs1$14$ , \picorv32_core/pcpi_rs2$14$ );  // ../src/picorv32.v(1230)
  AL_MUX \picorv32_core/u537  (
    .i0(\picorv32_core/mem_do_rinst ),
    .i1(\picorv32_core/mem_do_prefetch ),
    .sel(\picorv32_core/n553 ),
    .o(\picorv32_core/n568 ));  // ../src/picorv32.v(1789)
  not \picorv32_core/u538  (\picorv32_core/n572 , \picorv32_core/mem_do_prefetch );  // ../src/picorv32.v(1795)
  or \picorv32_core/u539  (\picorv32_core/n597 , \picorv32_core/n572 , \picorv32_core/mem_done );  // ../src/picorv32.v(1795)
  not \picorv32_core/u540  (\picorv32_core/n574 , \picorv32_core/mem_do_wdata );  // ../src/picorv32.v(1796)
  or \picorv32_core/u544  (\picorv32_core/n441 [13], \picorv32_core/pcpi_rs1$13$ , \picorv32_core/pcpi_rs2$13$ );  // ../src/picorv32.v(1230)
  and \picorv32_core/u545  (\picorv32_core/n580 , \picorv32_core/n572 , \picorv32_core/mem_done );  // ../src/picorv32.v(1810)
  and \picorv32_core/u548  (\picorv32_core/n443 [27], \picorv32_core/pcpi_rs1$27$ , \picorv32_core/pcpi_rs2$27$ );  // ../src/picorv32.v(1232)
  and \picorv32_core/u549  (\picorv32_core/n443 [28], \picorv32_core/pcpi_rs1$28$ , \picorv32_core/pcpi_rs2$28$ );  // ../src/picorv32.v(1232)
  and \picorv32_core/u550  (\picorv32_core/n443 [29], \picorv32_core/pcpi_rs1$29$ , \picorv32_core/pcpi_rs2$29$ );  // ../src/picorv32.v(1232)
  or \picorv32_core/u551  (\picorv32_core/n441 [12], \picorv32_core/pcpi_rs1$12$ , \picorv32_core/pcpi_rs2$12$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u552  (\picorv32_core/n441 [11], \picorv32_core/pcpi_rs1$11$ , \picorv32_core/pcpi_rs2$11$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u553  (\picorv32_core/n441 [10], \picorv32_core/pcpi_rs1$10$ , \picorv32_core/pcpi_rs2$10$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u554  (\picorv32_core/n599 , \picorv32_core/instr_lb , \picorv32_core/instr_lbu );  // ../src/picorv32.v(1824)
  or \picorv32_core/u555  (\picorv32_core/n600 , \picorv32_core/instr_lh , \picorv32_core/instr_lhu );  // ../src/picorv32.v(1825)
  or \picorv32_core/u559  (\picorv32_core/n441 [9], \picorv32_core/pcpi_rs1$9$ , \picorv32_core/pcpi_rs2$9$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u563  (\picorv32_core/n441 [8], \picorv32_core/pcpi_rs1$8$ , \picorv32_core/pcpi_rs2$8$ );  // ../src/picorv32.v(1230)
  or \picorv32_core/u564  (\picorv32_core/n441 [7], \picorv32_core/pcpi_rs1$7$ , mem_la_wdata[7]);  // ../src/picorv32.v(1230)
  or \picorv32_core/u568  (\picorv32_core/n441 [6], \picorv32_core/pcpi_rs1$6$ , mem_la_wdata[6]);  // ../src/picorv32.v(1230)
  or \picorv32_core/u569  (\picorv32_core/n441 [5], \picorv32_core/pcpi_rs1$5$ , mem_la_wdata[5]);  // ../src/picorv32.v(1230)
  not \picorv32_core/u57  (\picorv32_core/n135 [0], \picorv32_core/n10 );  // ../src/picorv32.v(581)
  and \picorv32_core/u570  (\picorv32_core/n443 [22], \picorv32_core/pcpi_rs1$22$ , \picorv32_core/pcpi_rs2$22$ );  // ../src/picorv32.v(1232)
  AL_MUX \picorv32_core/u571  (
    .i0(\picorv32_core/latched_is_lu ),
    .i1(\picorv32_core/is_lbu_lhu_lw ),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n653 ));
  AL_MUX \picorv32_core/u572  (
    .i0(\picorv32_core/latched_is_lh ),
    .i1(\picorv32_core/instr_lh ),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n654 ));
  AL_MUX \picorv32_core/u573  (
    .i0(\picorv32_core/latched_is_lb ),
    .i1(\picorv32_core/instr_lb ),
    .sel(\picorv32_core/mux132_b0_sel_is_3_o ),
    .o(\picorv32_core/n655 ));
  and \picorv32_core/u574  (\picorv32_core/n443 [23], \picorv32_core/pcpi_rs1$23$ , \picorv32_core/pcpi_rs2$23$ );  // ../src/picorv32.v(1232)
  AL_MUX \picorv32_core/u576  (
    .i0(\picorv32_core/n170 ),
    .i1(1'b1),
    .sel(\picorv32_core/mux148_b0_sel_is_3_o ),
    .o(\picorv32_core/n659 ));
  or \picorv32_core/u578  (\picorv32_core/n441 [4], \picorv32_core/pcpi_rs1$4$ , mem_la_wdata[4]);  // ../src/picorv32.v(1230)
  or \picorv32_core/u579  (\picorv32_core/n448 , \picorv32_core/is_rdcycle_rdcycleh_rdinstr_rdinstrh , \picorv32_core/instr_trap );  // ../src/picorv32.v(1694)
  or \picorv32_core/u580  (\picorv32_core/n684 , \picorv32_core/n669 , \picorv32_core/n668 );  // ../src/picorv32.v(1851)
  or \picorv32_core/u581  (\picorv32_core/n676 , \picorv32_core/n667 , \picorv32_core/n669 );  // ../src/picorv32.v(1851)
  or \picorv32_core/u582  (\picorv32_core/n686 , \picorv32_core/n665 , \picorv32_core/n662 );  // ../src/picorv32.v(1851)
  or \picorv32_core/u583  (\picorv32_core/n441 [3], \picorv32_core/pcpi_rs1$3$ , mem_la_wdata[3]);  // ../src/picorv32.v(1230)
  or \picorv32_core/u584  (\picorv32_core/n594 , \picorv32_core/n668 , \picorv32_core/n667 );  // ../src/picorv32.v(1851)
  or \picorv32_core/u585  (\picorv32_core/n441 [2], \picorv32_core/pcpi_rs1$2$ , mem_la_wdata[2]);  // ../src/picorv32.v(1230)
  or \picorv32_core/u586  (\picorv32_core/n441 [1], \picorv32_core/pcpi_rs1$1$ , mem_la_wdata[1]);  // ../src/picorv32.v(1230)
  and \picorv32_core/u589_sel_is_3  (\picorv32_core/u589_sel_is_3_o , \picorv32_core/n663 , \picorv32_core/mux127_b0_sel_is_1_o );
  not \picorv32_core/u59  (\picorv32_core/n353 , \picorv32_core/pcpi_rs1$0$ );  // ../src/picorv32.v(383)
  or \picorv32_core/u595  (\picorv32_core/n589 , \picorv32_core/n667 , \picorv32_core/n666 );  // ../src/picorv32.v(1851)
  and \picorv32_core/u596_sel_is_3  (\picorv32_core/u596_sel_is_3_o , \picorv32_core/n666 , \picorv32_core/is_beq_bne_blt_bge_bltu_bgeu );
  and \picorv32_core/u597_sel_is_3  (\picorv32_core/u597_sel_is_3_o , \picorv32_core/n668 , \picorv32_core/n597 );
  or \picorv32_core/u598  (\picorv32_core/n592 , \picorv32_core/n667 , \picorv32_core/n665 );  // ../src/picorv32.v(1851)
  and \picorv32_core/u599_sel_is_3  (\picorv32_core/u599_sel_is_3_o , \picorv32_core/n669 , \picorv32_core/n597 );
  not \picorv32_core/u60  (\picorv32_core/n21 , \picorv32_core/n8 );  // ../src/picorv32.v(343)
  and \picorv32_core/u61  (\picorv32_core/n43 , \picorv32_core/mem_done , \picorv32_core/n0 );  // ../src/picorv32.v(400)
  AL_MUX \picorv32_core/u615  (
    .i0(\picorv32_core/n671 ),
    .i1(\picorv32_core/mem_do_rinst ),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n718 ));  // ../src/picorv32.v(1851)
  and \picorv32_core/u616_sel_is_2  (\picorv32_core/u616_sel_is_2_o , resetn, \picorv32_core/n663 );
  and \picorv32_core/u617_sel_is_2  (\picorv32_core/u617_sel_is_2_o , resetn, \picorv32_core/u589_sel_is_3_o );
  and \picorv32_core/u62  (\picorv32_core/n443 [21], \picorv32_core/pcpi_rs1$21$ , \picorv32_core/pcpi_rs2$21$ );  // ../src/picorv32.v(1232)
  AL_MUX \picorv32_core/u622  (
    .i0(\picorv32_core/n698 ),
    .i1(\picorv32_core/n170 ),
    .sel(\picorv32_core/n407 ),
    .o(\picorv32_core/n727 ));  // ../src/picorv32.v(1851)
  AL_MUX \picorv32_core/u623  (
    .i0(1'b0),
    .i1(\picorv32_core/alu_out_0 ),
    .sel(\picorv32_core/u623_sel_is_2_o ),
    .o(\picorv32_core/n728 ));
  and \picorv32_core/u623_sel_is_2  (\picorv32_core/u623_sel_is_2_o , resetn, \picorv32_core/u596_sel_is_3_o );
  AL_MUX \picorv32_core/u624  (
    .i0(1'b0),
    .i1(\picorv32_core/n574 ),
    .sel(\picorv32_core/u624_sel_is_2_o ),
    .o(\picorv32_core/n729 ));
  and \picorv32_core/u624_sel_is_2  (\picorv32_core/u624_sel_is_2_o , resetn, \picorv32_core/u597_sel_is_3_o );
  and \picorv32_core/u625_sel_is_2  (\picorv32_core/u625_sel_is_2_o , resetn, \picorv32_core/sel46_sel_is_2_o );
  AL_MUX \picorv32_core/u626  (
    .i0(1'b0),
    .i1(\picorv32_core/n598 ),
    .sel(\picorv32_core/u626_sel_is_2_o ),
    .o(\picorv32_core/n731 ));
  and \picorv32_core/u626_sel_is_2  (\picorv32_core/u626_sel_is_2_o , resetn, \picorv32_core/u599_sel_is_3_o );
  or \picorv32_core/u627  (\picorv32_core/n732 , \picorv32_core/mem_do_rdata , \picorv32_core/mem_do_wdata );  // ../src/picorv32.v(1853)
  and \picorv32_core/u628  (\picorv32_core/n733 , resetn, \picorv32_core/n732 );  // ../src/picorv32.v(1853)
  and \picorv32_core/u629  (\picorv32_core/n736 , \picorv32_core/n734 , \picorv32_core/n735 );  // ../src/picorv32.v(1854)
  and \picorv32_core/u63  (\picorv32_core/n443 [25], \picorv32_core/pcpi_rs1$25$ , \picorv32_core/pcpi_rs2$25$ );  // ../src/picorv32.v(1232)
  and \picorv32_core/u630  (\picorv32_core/n740 , \picorv32_core/n738 , \picorv32_core/n739 );  // ../src/picorv32.v(1861)
  and \picorv32_core/u631  (\picorv32_core/n743 , resetn, \picorv32_core/mem_do_rinst );  // ../src/picorv32.v(1869)
  and \picorv32_core/u632  (\picorv32_core/n744 , \picorv32_core/n743 , \picorv32_core/reg_pc [0]);  // ../src/picorv32.v(1869)
  and \picorv32_core/u633  (\picorv32_core/n443 [31], \picorv32_core/pcpi_rs1$31$ , \picorv32_core/pcpi_rs2$31$ );  // ../src/picorv32.v(1232)
  or \picorv32_core/u634  (\picorv32_core/n747 , \picorv32_core/n407 , \picorv32_core/mem_done );  // ../src/picorv32.v(1880)
  AL_MUX \picorv32_core/u636  (
    .i0(\picorv32_core/n718 ),
    .i1(1'b0),
    .sel(\picorv32_core/n747 ),
    .o(\picorv32_core/n749 ));  // ../src/picorv32.v(1885)
  AL_MUX \picorv32_core/u64  (
    .i0(\picorv32_core/n353 ),
    .i1(1'b0),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n40 [0]));  // ../src/picorv32.v(383)
  or \picorv32_core/u65  (\picorv32_core/n701 , \picorv32_core/n46 , \picorv32_core/n593 );  // ../src/picorv32.v(1851)
  AL_MUX \picorv32_core/u66  (
    .i0(\picorv32_core/pcpi_rs1$0$ ),
    .i1(1'b0),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n40 [1]));  // ../src/picorv32.v(383)
  not \picorv32_core/u663  (\picorv32_core/n38 [0], \picorv32_core/pcpi_rs1$1$ );  // ../src/picorv32.v(375)
  and \picorv32_core/u664  (\picorv32_core/n443 [30], \picorv32_core/pcpi_rs1$30$ , \picorv32_core/pcpi_rs2$30$ );  // ../src/picorv32.v(1232)
  AL_MUX \picorv32_core/u68  (
    .i0(1'b0),
    .i1(\picorv32_core/n353 ),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n40 [2]));  // ../src/picorv32.v(383)
  and \picorv32_core/u7  (\picorv32_core/mem_la_firstword , \picorv32_core/n1 , \picorv32_core/mem_la_secondword_neg );  // ../src/picorv32.v(326)
  and \picorv32_core/u70  (\picorv32_core/n443 [26], \picorv32_core/pcpi_rs1$26$ , \picorv32_core/pcpi_rs2$26$ );  // ../src/picorv32.v(1232)
  or \picorv32_core/u71  (\picorv32_core/n50 , \picorv32_core/n99 , \picorv32_core/n44 );  // ../src/picorv32.v(416)
  AL_MUX \picorv32_core/u72  (
    .i0(1'b0),
    .i1(\picorv32_core/pcpi_rs1$0$ ),
    .sel(\picorv32_core/pcpi_rs1$1$ ),
    .o(\picorv32_core/n40 [3]));  // ../src/picorv32.v(383)
  and \picorv32_core/u73  (\picorv32_core/n443 [18], \picorv32_core/pcpi_rs1$18$ , \picorv32_core/pcpi_rs2$18$ );  // ../src/picorv32.v(1232)
  and \picorv32_core/u74  (\picorv32_core/n443 [19], \picorv32_core/pcpi_rs1$19$ , \picorv32_core/pcpi_rs2$19$ );  // ../src/picorv32.v(1232)
  and \picorv32_core/u75  (\picorv32_core/n443 [20], \picorv32_core/pcpi_rs1$20$ , \picorv32_core/pcpi_rs2$20$ );  // ../src/picorv32.v(1232)
  or \picorv32_core/u76  (\picorv32_core/n697 , \picorv32_core/n592 , \picorv32_core/n593 );  // ../src/picorv32.v(1851)
  and \picorv32_core/u79  (\picorv32_core/n74 , \picorv32_core/n72 , \picorv32_core/n73 );  // ../src/picorv32.v(483)
  or \picorv32_core/u80  (\picorv32_core/n633 , \picorv32_core/decoded_rs1 [2], \picorv32_core/n639 );  // ../src/picorv32.v(1328)
  or \picorv32_core/u81  (\picorv32_core/n457 , \picorv32_core/n640 , \picorv32_core/n633 );  // ../src/picorv32.v(1328)
  or \picorv32_core/u83  (\picorv32_core/n588 , \picorv32_core/n668 , \picorv32_core/n589 );  // ../src/picorv32.v(1851)
  or \picorv32_core/u86  (\picorv32_core/n682 , \picorv32_core/n588 , \picorv32_core/n746 );  // ../src/picorv32.v(1851)
  and \picorv32_core/u87  (\picorv32_core/n443 [1], \picorv32_core/pcpi_rs1$1$ , mem_la_wdata[1]);  // ../src/picorv32.v(1232)
  or \picorv32_core/u88  (\picorv32_core/n650 , \picorv32_core/is_jalr_addi_slti_sltiu_xori_ori_andi , \picorv32_core/n651 );  // ../src/picorv32.v(1694)
  and \picorv32_core/u91  (\picorv32_core/n80 , \picorv32_core/n72 , \picorv32_core/n79 );  // ../src/picorv32.v(487)
  and \picorv32_core/u92  (\picorv32_core/n443 [2], \picorv32_core/pcpi_rs1$2$ , mem_la_wdata[2]);  // ../src/picorv32.v(1232)
  and \picorv32_core/u93  (\picorv32_core/n443 [3], \picorv32_core/pcpi_rs1$3$ , mem_la_wdata[3]);  // ../src/picorv32.v(1232)
  and \picorv32_core/u94  (\picorv32_core/n443 [4], \picorv32_core/pcpi_rs1$4$ , mem_la_wdata[4]);  // ../src/picorv32.v(1232)
  and \picorv32_core/u95  (\picorv32_core/n443 [5], \picorv32_core/pcpi_rs1$5$ , mem_la_wdata[5]);  // ../src/picorv32.v(1232)
  or \picorv32_core/u96  (\picorv32_core/n648 , \picorv32_core/is_lui_auipc_jal , \picorv32_core/n448 );  // ../src/picorv32.v(1694)
  or \picorv32_core/u97  (\picorv32_core/n647 , \picorv32_core/n650 , \picorv32_core/n648 );  // ../src/picorv32.v(1694)
  and \picorv32_core/u98  (\picorv32_core/n86 , \picorv32_core/n84 , \picorv32_core/n85 );  // ../src/picorv32.v(491)
  reg_ar_as_w1 reg0_b0 (
    .clk(clk),
    .d(n3[0]),
    .en(n2),
    .reset(1'b0),
    .set(1'b0),
    .q(initial_reset[0]));  // ../src/top.v(42)
  reg_ar_as_w1 reg0_b1 (
    .clk(clk),
    .d(n3[1]),
    .en(n2),
    .reset(1'b0),
    .set(1'b0),
    .q(initial_reset[1]));  // ../src/top.v(42)
  reg_ar_as_w1 reg1_b0 (
    .clk(clk),
    .d(n17[0]),
    .en(n16),
    .reset(1'b0),
    .set(~resetn),
    .q(out_byte[0]));  // ../src/top.v(128)
  reg_ar_as_w1 reg1_b1 (
    .clk(clk),
    .d(n17[1]),
    .en(n16),
    .reset(1'b0),
    .set(~resetn),
    .q(out_byte[1]));  // ../src/top.v(128)
  reg_ar_as_w1 reg1_b2 (
    .clk(clk),
    .d(n17[2]),
    .en(n16),
    .reset(1'b0),
    .set(~resetn),
    .q(out_byte[2]));  // ../src/top.v(128)
  reg_ar_as_w1 reg1_b3 (
    .clk(clk),
    .d(n17[3]),
    .en(n16),
    .reset(1'b0),
    .set(~resetn),
    .q(out_byte[3]));  // ../src/top.v(128)
  reg_ar_as_w1 reg1_b4 (
    .clk(clk),
    .d(n17[4]),
    .en(n16),
    .reset(1'b0),
    .set(~resetn),
    .q(out_byte[4]));  // ../src/top.v(128)
  reg_ar_as_w1 reg1_b5 (
    .clk(clk),
    .d(n17[5]),
    .en(n16),
    .reset(1'b0),
    .set(~resetn),
    .q(out_byte[5]));  // ../src/top.v(128)
  reg_ar_as_w1 reg1_b6 (
    .clk(clk),
    .d(n17[6]),
    .en(n16),
    .reset(1'b0),
    .set(~resetn),
    .q(out_byte[6]));  // ../src/top.v(128)
  reg_ar_as_w1 reg1_b7 (
    .clk(clk),
    .d(n17[7]),
    .en(n16),
    .reset(1'b0),
    .set(~resetn),
    .q(out_byte[7]));  // ../src/top.v(128)
  reg_ar_as_w1 resetn_reg (
    .clk(clk),
    .d(n1),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(resetn));  // ../src/top.v(42)
  not u11 (n17[5], mem_la_wdata[5]);  // ../src/top.v(126)
  and u12 (n11, \picorv32_core/n116 [2], n6);  // ../src/top.v(88)
  not u13 (n17[4], mem_la_wdata[4]);  // ../src/top.v(126)
  not u15 (n17[3], mem_la_wdata[3]);  // ../src/top.v(126)
  and u16 (n13, \picorv32_core/n116 [3], n6);  // ../src/top.v(95)
  not u17 (n17[2], mem_la_wdata[2]);  // ../src/top.v(126)
  not u18 (n17[1], mem_la_wdata[1]);  // ../src/top.v(126)
  and u19 (n16, mem_la_write, n15);  // ../src/top.v(124)
  and u2 (n1, resetn_i, n0);  // ../src/top.v(38)
  not u20 (n17[0], mem_la_wdata[0]);  // ../src/top.v(126)
  and u4 (n7, \picorv32_core/n116 [0], n6);  // ../src/top.v(74)
  not u7 (n17[7], mem_la_wdata[7]);  // ../src/top.v(126)
  and u8 (n9, \picorv32_core/n116 [1], n6);  // ../src/top.v(81)
  not u9 (n17[6], mem_la_wdata[6]);  // ../src/top.v(126)
  add_pu32_pu32_o32 \uart/add0  (
    .i0(\uart/uart_counter ),
    .i1(32'b00000000000000000000000000000001),
    .o(\uart/n5 ));  // ../src/uart.v(68)
  add_pu4_pu4_o4 \uart/add1  (
    .i0(\uart/uart_status_txd ),
    .i1(4'b0001),
    .o(\uart/n35 ));  // ../src/uart.v(133)
  add_pu4_pu4_o4 \uart/add2  (
    .i0(\uart/uart_smp_rx ),
    .i1(4'b0001),
    .o(\uart/n49 ));  // ../src/uart.v(194)
  add_pu4_pu4_o4 \uart/add3  (
    .i0(\uart/uart_status_rxd ),
    .i1(4'b0001),
    .o(\uart/n77 ));  // ../src/uart.v(231)
  eq_w4 \uart/eq0  (
    .i0(\uart/uart_status_txd ),
    .i1(4'b0000),
    .o(\uart/n9 ));  // ../src/uart.v(80)
  eq_w3 \uart/eq1  (
    .i0(\uart/uart_cnt_rx ),
    .i1(3'b100),
    .o(\uart/n51 ));  // ../src/uart.v(197)
  eq_w3 \uart/eq2  (
    .i0(\uart/uart_cnt_rx ),
    .i1(3'b010),
    .o(\uart/n90 ));  // ../src/uart.v(241)
  lt_u32_u32 \uart/lt0  (
    .ci(1'b1),
    .i0(\uart/uart_bsrr ),
    .i1(\uart/uart_counter ),
    .o(\uart/n2 ));  // ../src/uart.v(59)
  lt_u4_u4 \uart/lt1  (
    .ci(1'b1),
    .i0(4'b0010),
    .i1(\uart/uart_smp_rx ),
    .o(\uart/n52 ));  // ../src/uart.v(200)
  binary_mux_s1_w1 \uart/mux0_b0  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\uart/n3 ),
    .o(\uart/n4 [0]));  // ../src/uart.v(63)
  binary_mux_s1_w1 \uart/mux0_b1  (
    .i0(1'b0),
    .i1(\uart/uart_op_clock_by_3_c [0]),
    .sel(\uart/n3 ),
    .o(\uart/n4 [1]));  // ../src/uart.v(63)
  and \uart/mux10_b0_sel_is_3  (\uart/mux10_b0_sel_is_3_o , mem_la_write, \uart/mux6_b0_sel_is_4_o );
  and \uart/mux12_b0_sel_is_3  (\uart/mux12_b0_sel_is_3_o , uart_sel, \uart/mux9_b0_sel_is_3_o );
  and \uart/mux13_b0_sel_is_3  (\uart/mux13_b0_sel_is_3_o , uart_sel, \uart/mux10_b0_sel_is_3_o );
  and \uart/mux14_b0_sel_is_1  (\uart/mux14_b0_sel_is_1_o , uart_sel, mem_la_write_neg);
  and \uart/mux15_b0_sel_is_2  (\uart/mux15_b0_sel_is_2_o , resetn, \uart/mux13_b0_sel_is_3_o );
  binary_mux_s3_w1 \uart/mux16  (
    .i0(\uart/uart_odr [0]),
    .i1(\uart/uart_odr [1]),
    .i2(\uart/uart_odr [2]),
    .i3(\uart/uart_odr [3]),
    .i4(\uart/uart_odr [4]),
    .i5(\uart/uart_odr [5]),
    .i6(\uart/uart_odr [6]),
    .i7(\uart/uart_odr [7]),
    .sel(\uart/n33 [2:0]),
    .o(\uart/n34 ));  // ../src/uart.v(131)
  binary_mux_s4_w1 \uart/mux17_b0  (
    .i0(\uart/n31 [0]),
    .i1(\uart/n37 [0]),
    .i10(\uart/n37 [0]),
    .i11(1'b0),
    .i12(1'b0),
    .i13(1'b0),
    .i14(1'b0),
    .i15(1'b0),
    .i2(\uart/n36 [0]),
    .i3(\uart/n36 [0]),
    .i4(\uart/n36 [0]),
    .i5(\uart/n36 [0]),
    .i6(\uart/n36 [0]),
    .i7(\uart/n36 [0]),
    .i8(\uart/n36 [0]),
    .i9(\uart/n36 [0]),
    .sel(\uart/uart_status_txd ),
    .o(\uart/n38 [0]));  // ../src/uart.v(143)
  binary_mux_s4_w1 \uart/mux17_b1  (
    .i0(\uart/n31 [1]),
    .i1(\uart/n32 [1]),
    .i10(\uart/n31 [1]),
    .i11(1'b0),
    .i12(1'b0),
    .i13(1'b0),
    .i14(1'b0),
    .i15(1'b0),
    .i2(\uart/n36 [1]),
    .i3(\uart/n36 [1]),
    .i4(\uart/n36 [1]),
    .i5(\uart/n36 [1]),
    .i6(\uart/n36 [1]),
    .i7(\uart/n36 [1]),
    .i8(\uart/n36 [1]),
    .i9(\uart/n36 [1]),
    .sel(\uart/uart_status_txd ),
    .o(\uart/n38 [1]));  // ../src/uart.v(143)
  binary_mux_s4_w1 \uart/mux17_b2  (
    .i0(\uart/n37 [2]),
    .i1(\uart/n37 [2]),
    .i10(\uart/n37 [2]),
    .i11(1'b0),
    .i12(1'b0),
    .i13(1'b0),
    .i14(1'b0),
    .i15(1'b0),
    .i2(\uart/n36 [2]),
    .i3(\uart/n36 [2]),
    .i4(\uart/n36 [2]),
    .i5(\uart/n36 [2]),
    .i6(\uart/n36 [2]),
    .i7(\uart/n36 [2]),
    .i8(\uart/n36 [2]),
    .i9(\uart/n36 [2]),
    .sel(\uart/uart_status_txd ),
    .o(\uart/n38 [2]));  // ../src/uart.v(143)
  binary_mux_s4_w1 \uart/mux17_b3  (
    .i0(\uart/n37 [3]),
    .i1(\uart/n37 [3]),
    .i10(\uart/n37 [3]),
    .i11(1'b0),
    .i12(1'b0),
    .i13(1'b0),
    .i14(1'b0),
    .i15(1'b0),
    .i2(\uart/n36 [3]),
    .i3(\uart/n36 [3]),
    .i4(\uart/n36 [3]),
    .i5(\uart/n36 [3]),
    .i6(\uart/n36 [3]),
    .i7(\uart/n36 [3]),
    .i8(\uart/n36 [3]),
    .i9(\uart/n36 [3]),
    .sel(\uart/uart_status_txd ),
    .o(\uart/n38 [3]));  // ../src/uart.v(143)
  binary_mux_s4_w1 \uart/mux18  (
    .i0(txd),
    .i1(1'b0),
    .i10(1'b1),
    .i11(txd),
    .i12(txd),
    .i13(txd),
    .i14(txd),
    .i15(txd),
    .i2(\uart/n34 ),
    .i3(\uart/n34 ),
    .i4(\uart/n34 ),
    .i5(\uart/n34 ),
    .i6(\uart/n34 ),
    .i7(\uart/n34 ),
    .i8(\uart/n34 ),
    .i9(\uart/n34 ),
    .sel(\uart/uart_status_txd ),
    .o(\uart/n39 ));  // ../src/uart.v(143)
  binary_mux_s1_w1 \uart/mux1_b0  (
    .i0(\uart/n5 [0]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [0]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b1  (
    .i0(\uart/n5 [1]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [1]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b10  (
    .i0(\uart/n5 [10]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [10]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b11  (
    .i0(\uart/n5 [11]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [11]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b12  (
    .i0(\uart/n5 [12]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [12]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b13  (
    .i0(\uart/n5 [13]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [13]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b14  (
    .i0(\uart/n5 [14]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [14]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b15  (
    .i0(\uart/n5 [15]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [15]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b16  (
    .i0(\uart/n5 [16]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [16]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b17  (
    .i0(\uart/n5 [17]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [17]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b18  (
    .i0(\uart/n5 [18]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [18]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b19  (
    .i0(\uart/n5 [19]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [19]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b2  (
    .i0(\uart/n5 [2]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [2]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b20  (
    .i0(\uart/n5 [20]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [20]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b21  (
    .i0(\uart/n5 [21]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [21]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b22  (
    .i0(\uart/n5 [22]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [22]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b23  (
    .i0(\uart/n5 [23]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [23]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b24  (
    .i0(\uart/n5 [24]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [24]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b25  (
    .i0(\uart/n5 [25]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [25]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b26  (
    .i0(\uart/n5 [26]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [26]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b27  (
    .i0(\uart/n5 [27]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [27]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b28  (
    .i0(\uart/n5 [28]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [28]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b29  (
    .i0(\uart/n5 [29]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [29]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b3  (
    .i0(\uart/n5 [3]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [3]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b30  (
    .i0(\uart/n5 [30]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [30]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b31  (
    .i0(\uart/n5 [31]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [31]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b4  (
    .i0(\uart/n5 [4]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [4]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b5  (
    .i0(\uart/n5 [5]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [5]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b6  (
    .i0(\uart/n5 [6]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [6]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b7  (
    .i0(\uart/n5 [7]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [7]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b8  (
    .i0(\uart/n5 [8]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [8]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux1_b9  (
    .i0(\uart/n5 [9]),
    .i1(1'b0),
    .sel(\uart/n2 ),
    .o(\uart/n6 [9]));  // ../src/uart.v(69)
  binary_mux_s1_w1 \uart/mux20_b0  (
    .i0(\uart/uart_idr_t [0]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n45 [0]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux20_b1  (
    .i0(\uart/uart_idr_t [1]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n45 [1]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux20_b2  (
    .i0(\uart/uart_idr_t [2]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n45 [2]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux20_b3  (
    .i0(\uart/uart_idr_t [3]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n45 [3]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux20_b4  (
    .i0(\uart/uart_idr_t [4]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n45 [4]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux20_b5  (
    .i0(\uart/uart_idr_t [5]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n45 [5]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux20_b6  (
    .i0(\uart/uart_idr_t [6]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n45 [6]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux20_b7  (
    .i0(\uart/uart_idr_t [7]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n45 [7]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux21_b0  (
    .i0(\uart/uart_cnt_rx [0]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n46 [0]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux21_b1  (
    .i0(\uart/uart_cnt_rx [1]),
    .i1(1'b1),
    .sel(\uart/n44 ),
    .o(\uart/n46 [1]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux21_b2  (
    .i0(\uart/uart_cnt_rx [2]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n46 [2]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux22_b0  (
    .i0(\uart/uart_smp_rx [0]),
    .i1(1'b1),
    .sel(\uart/n44 ),
    .o(\uart/n47 [0]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux22_b1  (
    .i0(\uart/uart_smp_rx [1]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n47 [1]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux22_b2  (
    .i0(\uart/uart_smp_rx [2]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n47 [2]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux22_b3  (
    .i0(\uart/uart_smp_rx [3]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n47 [3]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux23_b0  (
    .i0(\uart/uart_status_rxd [0]),
    .i1(1'b1),
    .sel(\uart/n44 ),
    .o(\uart/n48 [0]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux23_b1  (
    .i0(\uart/uart_status_rxd [1]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n48 [1]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux23_b2  (
    .i0(\uart/uart_status_rxd [2]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n48 [2]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux23_b3  (
    .i0(\uart/uart_status_rxd [3]),
    .i1(1'b0),
    .sel(\uart/n44 ),
    .o(\uart/n48 [3]));  // ../src/uart.v(188)
  binary_mux_s1_w1 \uart/mux24_b0  (
    .i0(\uart/n49 [0]),
    .i1(\uart/uart_smp_rx [0]),
    .sel(rxd),
    .o(\uart/n50 [0]));  // ../src/uart.v(195)
  binary_mux_s1_w1 \uart/mux24_b1  (
    .i0(\uart/n49 [1]),
    .i1(\uart/uart_smp_rx [1]),
    .sel(rxd),
    .o(\uart/n50 [1]));  // ../src/uart.v(195)
  binary_mux_s1_w1 \uart/mux24_b2  (
    .i0(\uart/n49 [2]),
    .i1(\uart/uart_smp_rx [2]),
    .sel(rxd),
    .o(\uart/n50 [2]));  // ../src/uart.v(195)
  binary_mux_s1_w1 \uart/mux24_b3  (
    .i0(\uart/n49 [3]),
    .i1(\uart/uart_smp_rx [3]),
    .sel(rxd),
    .o(\uart/n50 [3]));  // ../src/uart.v(195)
  binary_mux_s1_w1 \uart/mux26_b0  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\uart/n56 ),
    .o(\uart/n81 [0]));  // ../src/uart.v(209)
  binary_mux_s1_w1 \uart/mux26_b1  (
    .i0(1'b0),
    .i1(\uart/uart_cnt_rx [0]),
    .sel(\uart/n56 ),
    .o(\uart/n81 [1]));  // ../src/uart.v(209)
  binary_mux_s1_w1 \uart/mux26_b2  (
    .i0(1'b0),
    .i1(\uart/uart_cnt_rx [1]),
    .sel(\uart/n56 ),
    .o(\uart/n81 [2]));  // ../src/uart.v(209)
  binary_mux_s1_w1 \uart/mux27_b0  (
    .i0(\uart/uart_idr_t [6]),
    .i1(1'b0),
    .sel(\uart/n62 ),
    .o(\uart/n63 [0]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux27_b1  (
    .i0(\uart/uart_idr_t [6]),
    .i1(1'b1),
    .sel(\uart/n62 ),
    .o(\uart/n63 [1]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux28_b0  (
    .i0(\uart/uart_idr_t [5]),
    .i1(1'b0),
    .sel(\uart/n64 ),
    .o(\uart/n65 [0]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux28_b1  (
    .i0(\uart/uart_idr_t [5]),
    .i1(1'b1),
    .sel(\uart/n64 ),
    .o(\uart/n65 [1]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux29_b0  (
    .i0(\uart/uart_idr_t [4]),
    .i1(1'b0),
    .sel(\uart/n66 ),
    .o(\uart/n67 [0]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux29_b1  (
    .i0(\uart/uart_idr_t [4]),
    .i1(1'b1),
    .sel(\uart/n66 ),
    .o(\uart/n67 [1]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux30_b0  (
    .i0(\uart/uart_idr_t [3]),
    .i1(1'b0),
    .sel(\uart/n68 ),
    .o(\uart/n69 [0]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux30_b1  (
    .i0(\uart/uart_idr_t [3]),
    .i1(1'b1),
    .sel(\uart/n68 ),
    .o(\uart/n69 [1]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux31_b0  (
    .i0(\uart/uart_idr_t [2]),
    .i1(1'b0),
    .sel(\uart/n70 ),
    .o(\uart/n71 [0]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux31_b1  (
    .i0(\uart/uart_idr_t [2]),
    .i1(1'b1),
    .sel(\uart/n70 ),
    .o(\uart/n71 [1]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux32_b0  (
    .i0(\uart/uart_idr_t [1]),
    .i1(1'b0),
    .sel(\uart/n72 ),
    .o(\uart/n73 [0]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux32_b1  (
    .i0(\uart/uart_idr_t [1]),
    .i1(1'b1),
    .sel(\uart/n72 ),
    .o(\uart/n73 [1]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux33_b0  (
    .i0(\uart/uart_idr_t [0]),
    .i1(1'b0),
    .sel(\uart/n74 ),
    .o(\uart/n75 [0]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux33_b1  (
    .i0(\uart/uart_idr_t [0]),
    .i1(1'b1),
    .sel(\uart/n74 ),
    .o(\uart/n75 [1]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux34_b0  (
    .i0(\uart/n75 [1]),
    .i1(\uart/n75 [0]),
    .sel(\uart/n52 ),
    .o(\uart/n76 [0]));  // ../src/uart.v(229)
  binary_mux_s1_w1 \uart/mux34_b1  (
    .i0(\uart/n73 [1]),
    .i1(\uart/n73 [0]),
    .sel(\uart/n52 ),
    .o(\uart/n76 [1]));  // ../src/uart.v(229)
  binary_mux_s1_w1 \uart/mux34_b2  (
    .i0(\uart/n71 [1]),
    .i1(\uart/n71 [0]),
    .sel(\uart/n52 ),
    .o(\uart/n76 [2]));  // ../src/uart.v(229)
  binary_mux_s1_w1 \uart/mux34_b3  (
    .i0(\uart/n69 [1]),
    .i1(\uart/n69 [0]),
    .sel(\uart/n52 ),
    .o(\uart/n76 [3]));  // ../src/uart.v(229)
  binary_mux_s1_w1 \uart/mux34_b4  (
    .i0(\uart/n67 [1]),
    .i1(\uart/n67 [0]),
    .sel(\uart/n52 ),
    .o(\uart/n76 [4]));  // ../src/uart.v(229)
  binary_mux_s1_w1 \uart/mux34_b5  (
    .i0(\uart/n65 [1]),
    .i1(\uart/n65 [0]),
    .sel(\uart/n52 ),
    .o(\uart/n76 [5]));  // ../src/uart.v(229)
  binary_mux_s1_w1 \uart/mux34_b6  (
    .i0(\uart/n63 [1]),
    .i1(\uart/n63 [0]),
    .sel(\uart/n52 ),
    .o(\uart/n76 [6]));  // ../src/uart.v(229)
  binary_mux_s1_w1 \uart/mux34_b7  (
    .i0(\uart/n61 [1]),
    .i1(\uart/n61 [0]),
    .sel(\uart/n52 ),
    .o(\uart/n76 [7]));  // ../src/uart.v(229)
  binary_mux_s1_w1 \uart/mux35_b0  (
    .i0(\uart/uart_idr_t [0]),
    .i1(\uart/n76 [0]),
    .sel(\uart/n51 ),
    .o(\uart/n78 [0]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux35_b1  (
    .i0(\uart/uart_idr_t [1]),
    .i1(\uart/n76 [1]),
    .sel(\uart/n51 ),
    .o(\uart/n78 [1]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux35_b2  (
    .i0(\uart/uart_idr_t [2]),
    .i1(\uart/n76 [2]),
    .sel(\uart/n51 ),
    .o(\uart/n78 [2]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux35_b3  (
    .i0(\uart/uart_idr_t [3]),
    .i1(\uart/n76 [3]),
    .sel(\uart/n51 ),
    .o(\uart/n78 [3]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux35_b4  (
    .i0(\uart/uart_idr_t [4]),
    .i1(\uart/n76 [4]),
    .sel(\uart/n51 ),
    .o(\uart/n78 [4]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux35_b5  (
    .i0(\uart/uart_idr_t [5]),
    .i1(\uart/n76 [5]),
    .sel(\uart/n51 ),
    .o(\uart/n78 [5]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux35_b6  (
    .i0(\uart/uart_idr_t [6]),
    .i1(\uart/n76 [6]),
    .sel(\uart/n51 ),
    .o(\uart/n78 [6]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux35_b7  (
    .i0(\uart/uart_idr_t [7]),
    .i1(\uart/n76 [7]),
    .sel(\uart/n51 ),
    .o(\uart/n78 [7]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux36_b0  (
    .i0(\uart/uart_idr_t [7]),
    .i1(1'b0),
    .sel(\uart/n60 ),
    .o(\uart/n61 [0]));  // ../src/uart.v(227)
  binary_mux_s1_w1 \uart/mux36_b1  (
    .i0(\uart/uart_idr_t [7]),
    .i1(1'b1),
    .sel(\uart/n60 ),
    .o(\uart/n61 [1]));  // ../src/uart.v(227)
  AL_MUX \uart/mux37_b0  (
    .i0(\uart/n50 [0]),
    .i1(\uart/n44 ),
    .sel(\uart/mux37_b0_sel_is_3_o ),
    .o(\uart/n55 [0]));
  and \uart/mux37_b0_sel_is_3  (\uart/mux37_b0_sel_is_3_o , \uart/n51 , \uart/n52 );
  AL_MUX \uart/mux37_b1  (
    .i0(\uart/n50 [1]),
    .i1(1'b0),
    .sel(\uart/mux37_b0_sel_is_3_o ),
    .o(\uart/n55 [1]));
  AL_MUX \uart/mux37_b2  (
    .i0(\uart/n50 [2]),
    .i1(1'b0),
    .sel(\uart/mux37_b0_sel_is_3_o ),
    .o(\uart/n55 [2]));
  AL_MUX \uart/mux37_b3  (
    .i0(\uart/n50 [3]),
    .i1(1'b0),
    .sel(\uart/mux37_b0_sel_is_3_o ),
    .o(\uart/n55 [3]));
  binary_mux_s1_w1 \uart/mux37_b4  (
    .i0(\uart/n50 [0]),
    .i1(\uart/n44 ),
    .sel(\uart/n51 ),
    .o(\uart/n79 [0]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux37_b5  (
    .i0(\uart/n50 [1]),
    .i1(1'b0),
    .sel(\uart/n51 ),
    .o(\uart/n79 [1]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux37_b6  (
    .i0(\uart/n50 [2]),
    .i1(1'b0),
    .sel(\uart/n51 ),
    .o(\uart/n79 [2]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux37_b7  (
    .i0(\uart/n50 [3]),
    .i1(1'b0),
    .sel(\uart/n51 ),
    .o(\uart/n79 [3]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux38_b0  (
    .i0(\uart/uart_status_rxd [0]),
    .i1(1'b0),
    .sel(\uart/n90 ),
    .o(\uart/n92 [0]));  // ../src/uart.v(256)
  binary_mux_s1_w1 \uart/mux38_b1  (
    .i0(\uart/uart_status_rxd [1]),
    .i1(1'b0),
    .sel(\uart/n90 ),
    .o(\uart/n92 [1]));  // ../src/uart.v(256)
  binary_mux_s1_w1 \uart/mux38_b2  (
    .i0(\uart/uart_status_rxd [2]),
    .i1(1'b0),
    .sel(\uart/n90 ),
    .o(\uart/n92 [2]));  // ../src/uart.v(256)
  binary_mux_s1_w1 \uart/mux38_b3  (
    .i0(\uart/uart_status_rxd [3]),
    .i1(1'b0),
    .sel(\uart/n90 ),
    .o(\uart/n92 [3]));  // ../src/uart.v(256)
  binary_mux_s1_w1 \uart/mux40_b0  (
    .i0(\uart/uart_status_rxd [0]),
    .i1(1'b0),
    .sel(\uart/n51 ),
    .o(\uart/n54 [0]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux40_b1  (
    .i0(\uart/uart_status_rxd [1]),
    .i1(\uart/n52 ),
    .sel(\uart/n51 ),
    .o(\uart/n54 [1]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux40_b2  (
    .i0(\uart/uart_status_rxd [2]),
    .i1(1'b0),
    .sel(\uart/n51 ),
    .o(\uart/n54 [2]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux40_b3  (
    .i0(\uart/uart_status_rxd [3]),
    .i1(1'b0),
    .sel(\uart/n51 ),
    .o(\uart/n54 [3]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux40_b4  (
    .i0(\uart/uart_status_rxd [0]),
    .i1(\uart/n77 [0]),
    .sel(\uart/n51 ),
    .o(\uart/n80 [0]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux40_b5  (
    .i0(\uart/uart_status_rxd [1]),
    .i1(\uart/n77 [1]),
    .sel(\uart/n51 ),
    .o(\uart/n80 [1]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux40_b6  (
    .i0(\uart/uart_status_rxd [2]),
    .i1(\uart/n77 [2]),
    .sel(\uart/n51 ),
    .o(\uart/n80 [2]));  // ../src/uart.v(232)
  binary_mux_s1_w1 \uart/mux40_b7  (
    .i0(\uart/uart_status_rxd [3]),
    .i1(\uart/n77 [3]),
    .sel(\uart/n51 ),
    .o(\uart/n80 [3]));  // ../src/uart.v(232)
  binary_mux_s4_w1 \uart/mux41_b0  (
    .i0(\uart/n48 [0]),
    .i1(\uart/n54 [0]),
    .i10(\uart/n92 [0]),
    .i11(1'b0),
    .i12(1'b0),
    .i13(1'b0),
    .i14(1'b0),
    .i15(1'b0),
    .i2(\uart/n80 [0]),
    .i3(\uart/n80 [0]),
    .i4(\uart/n80 [0]),
    .i5(\uart/n80 [0]),
    .i6(\uart/n80 [0]),
    .i7(\uart/n80 [0]),
    .i8(\uart/n80 [0]),
    .i9(\uart/n80 [0]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n100 [0]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux41_b1  (
    .i0(\uart/n48 [1]),
    .i1(\uart/n54 [1]),
    .i10(\uart/n92 [1]),
    .i11(1'b0),
    .i12(1'b0),
    .i13(1'b0),
    .i14(1'b0),
    .i15(1'b0),
    .i2(\uart/n80 [1]),
    .i3(\uart/n80 [1]),
    .i4(\uart/n80 [1]),
    .i5(\uart/n80 [1]),
    .i6(\uart/n80 [1]),
    .i7(\uart/n80 [1]),
    .i8(\uart/n80 [1]),
    .i9(\uart/n80 [1]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n100 [1]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux41_b2  (
    .i0(\uart/n48 [2]),
    .i1(\uart/n54 [2]),
    .i10(\uart/n92 [2]),
    .i11(1'b0),
    .i12(1'b0),
    .i13(1'b0),
    .i14(1'b0),
    .i15(1'b0),
    .i2(\uart/n80 [2]),
    .i3(\uart/n80 [2]),
    .i4(\uart/n80 [2]),
    .i5(\uart/n80 [2]),
    .i6(\uart/n80 [2]),
    .i7(\uart/n80 [2]),
    .i8(\uart/n80 [2]),
    .i9(\uart/n80 [2]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n100 [2]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux41_b3  (
    .i0(\uart/n48 [3]),
    .i1(\uart/n54 [3]),
    .i10(\uart/n92 [3]),
    .i11(1'b0),
    .i12(1'b0),
    .i13(1'b0),
    .i14(1'b0),
    .i15(1'b0),
    .i2(\uart/n80 [3]),
    .i3(\uart/n80 [3]),
    .i4(\uart/n80 [3]),
    .i5(\uart/n80 [3]),
    .i6(\uart/n80 [3]),
    .i7(\uart/n80 [3]),
    .i8(\uart/n80 [3]),
    .i9(\uart/n80 [3]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n100 [3]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux42_b0  (
    .i0(\uart/n47 [0]),
    .i1(\uart/n55 [0]),
    .i10(\uart/n50 [0]),
    .i11(\uart/uart_smp_rx [0]),
    .i12(\uart/uart_smp_rx [0]),
    .i13(\uart/uart_smp_rx [0]),
    .i14(\uart/uart_smp_rx [0]),
    .i15(\uart/uart_smp_rx [0]),
    .i2(\uart/n79 [0]),
    .i3(\uart/n79 [0]),
    .i4(\uart/n79 [0]),
    .i5(\uart/n79 [0]),
    .i6(\uart/n79 [0]),
    .i7(\uart/n79 [0]),
    .i8(\uart/n79 [0]),
    .i9(\uart/n79 [0]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n101 [0]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux42_b1  (
    .i0(\uart/n47 [1]),
    .i1(\uart/n55 [1]),
    .i10(\uart/n50 [1]),
    .i11(\uart/uart_smp_rx [1]),
    .i12(\uart/uart_smp_rx [1]),
    .i13(\uart/uart_smp_rx [1]),
    .i14(\uart/uart_smp_rx [1]),
    .i15(\uart/uart_smp_rx [1]),
    .i2(\uart/n79 [1]),
    .i3(\uart/n79 [1]),
    .i4(\uart/n79 [1]),
    .i5(\uart/n79 [1]),
    .i6(\uart/n79 [1]),
    .i7(\uart/n79 [1]),
    .i8(\uart/n79 [1]),
    .i9(\uart/n79 [1]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n101 [1]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux42_b2  (
    .i0(\uart/n47 [2]),
    .i1(\uart/n55 [2]),
    .i10(\uart/n50 [2]),
    .i11(\uart/uart_smp_rx [2]),
    .i12(\uart/uart_smp_rx [2]),
    .i13(\uart/uart_smp_rx [2]),
    .i14(\uart/uart_smp_rx [2]),
    .i15(\uart/uart_smp_rx [2]),
    .i2(\uart/n79 [2]),
    .i3(\uart/n79 [2]),
    .i4(\uart/n79 [2]),
    .i5(\uart/n79 [2]),
    .i6(\uart/n79 [2]),
    .i7(\uart/n79 [2]),
    .i8(\uart/n79 [2]),
    .i9(\uart/n79 [2]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n101 [2]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux42_b3  (
    .i0(\uart/n47 [3]),
    .i1(\uart/n55 [3]),
    .i10(\uart/n50 [3]),
    .i11(\uart/uart_smp_rx [3]),
    .i12(\uart/uart_smp_rx [3]),
    .i13(\uart/uart_smp_rx [3]),
    .i14(\uart/uart_smp_rx [3]),
    .i15(\uart/uart_smp_rx [3]),
    .i2(\uart/n79 [3]),
    .i3(\uart/n79 [3]),
    .i4(\uart/n79 [3]),
    .i5(\uart/n79 [3]),
    .i6(\uart/n79 [3]),
    .i7(\uart/n79 [3]),
    .i8(\uart/n79 [3]),
    .i9(\uart/n79 [3]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n101 [3]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux43_b0  (
    .i0(\uart/n46 [0]),
    .i1(\uart/n81 [0]),
    .i10(\uart/n81 [0]),
    .i11(\uart/uart_cnt_rx [0]),
    .i12(\uart/uart_cnt_rx [0]),
    .i13(\uart/uart_cnt_rx [0]),
    .i14(\uart/uart_cnt_rx [0]),
    .i15(\uart/uart_cnt_rx [0]),
    .i2(\uart/n81 [0]),
    .i3(\uart/n81 [0]),
    .i4(\uart/n81 [0]),
    .i5(\uart/n81 [0]),
    .i6(\uart/n81 [0]),
    .i7(\uart/n81 [0]),
    .i8(\uart/n81 [0]),
    .i9(\uart/n81 [0]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n102 [0]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux43_b1  (
    .i0(\uart/n46 [1]),
    .i1(\uart/n81 [1]),
    .i10(\uart/n81 [1]),
    .i11(\uart/uart_cnt_rx [1]),
    .i12(\uart/uart_cnt_rx [1]),
    .i13(\uart/uart_cnt_rx [1]),
    .i14(\uart/uart_cnt_rx [1]),
    .i15(\uart/uart_cnt_rx [1]),
    .i2(\uart/n81 [1]),
    .i3(\uart/n81 [1]),
    .i4(\uart/n81 [1]),
    .i5(\uart/n81 [1]),
    .i6(\uart/n81 [1]),
    .i7(\uart/n81 [1]),
    .i8(\uart/n81 [1]),
    .i9(\uart/n81 [1]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n102 [1]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux43_b2  (
    .i0(\uart/n46 [2]),
    .i1(\uart/n81 [2]),
    .i10(\uart/n81 [2]),
    .i11(\uart/uart_cnt_rx [2]),
    .i12(\uart/uart_cnt_rx [2]),
    .i13(\uart/uart_cnt_rx [2]),
    .i14(\uart/uart_cnt_rx [2]),
    .i15(\uart/uart_cnt_rx [2]),
    .i2(\uart/n81 [2]),
    .i3(\uart/n81 [2]),
    .i4(\uart/n81 [2]),
    .i5(\uart/n81 [2]),
    .i6(\uart/n81 [2]),
    .i7(\uart/n81 [2]),
    .i8(\uart/n81 [2]),
    .i9(\uart/n81 [2]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n102 [2]));  // ../src/uart.v(261)
  and \uart/mux44_b0_sel_is_26  (\uart/mux44_b0_sel_is_26_o , \uart/uart_status_rxd$0$_neg , \uart/uart_status_rxd [1], \uart/uart_status_rxd$2$_neg , \uart/uart_status_rxd [3], \uart/n90 );
  binary_mux_s4_w1 \uart/mux47_b0  (
    .i0(\uart/n45 [0]),
    .i1(\uart/uart_idr_t [0]),
    .i10(\uart/uart_idr_t [0]),
    .i11(\uart/uart_idr_t [0]),
    .i12(\uart/uart_idr_t [0]),
    .i13(\uart/uart_idr_t [0]),
    .i14(\uart/uart_idr_t [0]),
    .i15(\uart/uart_idr_t [0]),
    .i2(\uart/n78 [0]),
    .i3(\uart/n78 [0]),
    .i4(\uart/n78 [0]),
    .i5(\uart/n78 [0]),
    .i6(\uart/n78 [0]),
    .i7(\uart/n78 [0]),
    .i8(\uart/n78 [0]),
    .i9(\uart/n78 [0]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n106 [0]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux47_b1  (
    .i0(\uart/n45 [1]),
    .i1(\uart/uart_idr_t [1]),
    .i10(\uart/uart_idr_t [1]),
    .i11(\uart/uart_idr_t [1]),
    .i12(\uart/uart_idr_t [1]),
    .i13(\uart/uart_idr_t [1]),
    .i14(\uart/uart_idr_t [1]),
    .i15(\uart/uart_idr_t [1]),
    .i2(\uart/n78 [1]),
    .i3(\uart/n78 [1]),
    .i4(\uart/n78 [1]),
    .i5(\uart/n78 [1]),
    .i6(\uart/n78 [1]),
    .i7(\uart/n78 [1]),
    .i8(\uart/n78 [1]),
    .i9(\uart/n78 [1]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n106 [1]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux47_b2  (
    .i0(\uart/n45 [2]),
    .i1(\uart/uart_idr_t [2]),
    .i10(\uart/uart_idr_t [2]),
    .i11(\uart/uart_idr_t [2]),
    .i12(\uart/uart_idr_t [2]),
    .i13(\uart/uart_idr_t [2]),
    .i14(\uart/uart_idr_t [2]),
    .i15(\uart/uart_idr_t [2]),
    .i2(\uart/n78 [2]),
    .i3(\uart/n78 [2]),
    .i4(\uart/n78 [2]),
    .i5(\uart/n78 [2]),
    .i6(\uart/n78 [2]),
    .i7(\uart/n78 [2]),
    .i8(\uart/n78 [2]),
    .i9(\uart/n78 [2]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n106 [2]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux47_b3  (
    .i0(\uart/n45 [3]),
    .i1(\uart/uart_idr_t [3]),
    .i10(\uart/uart_idr_t [3]),
    .i11(\uart/uart_idr_t [3]),
    .i12(\uart/uart_idr_t [3]),
    .i13(\uart/uart_idr_t [3]),
    .i14(\uart/uart_idr_t [3]),
    .i15(\uart/uart_idr_t [3]),
    .i2(\uart/n78 [3]),
    .i3(\uart/n78 [3]),
    .i4(\uart/n78 [3]),
    .i5(\uart/n78 [3]),
    .i6(\uart/n78 [3]),
    .i7(\uart/n78 [3]),
    .i8(\uart/n78 [3]),
    .i9(\uart/n78 [3]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n106 [3]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux47_b4  (
    .i0(\uart/n45 [4]),
    .i1(\uart/uart_idr_t [4]),
    .i10(\uart/uart_idr_t [4]),
    .i11(\uart/uart_idr_t [4]),
    .i12(\uart/uart_idr_t [4]),
    .i13(\uart/uart_idr_t [4]),
    .i14(\uart/uart_idr_t [4]),
    .i15(\uart/uart_idr_t [4]),
    .i2(\uart/n78 [4]),
    .i3(\uart/n78 [4]),
    .i4(\uart/n78 [4]),
    .i5(\uart/n78 [4]),
    .i6(\uart/n78 [4]),
    .i7(\uart/n78 [4]),
    .i8(\uart/n78 [4]),
    .i9(\uart/n78 [4]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n106 [4]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux47_b5  (
    .i0(\uart/n45 [5]),
    .i1(\uart/uart_idr_t [5]),
    .i10(\uart/uart_idr_t [5]),
    .i11(\uart/uart_idr_t [5]),
    .i12(\uart/uart_idr_t [5]),
    .i13(\uart/uart_idr_t [5]),
    .i14(\uart/uart_idr_t [5]),
    .i15(\uart/uart_idr_t [5]),
    .i2(\uart/n78 [5]),
    .i3(\uart/n78 [5]),
    .i4(\uart/n78 [5]),
    .i5(\uart/n78 [5]),
    .i6(\uart/n78 [5]),
    .i7(\uart/n78 [5]),
    .i8(\uart/n78 [5]),
    .i9(\uart/n78 [5]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n106 [5]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux47_b6  (
    .i0(\uart/n45 [6]),
    .i1(\uart/uart_idr_t [6]),
    .i10(\uart/uart_idr_t [6]),
    .i11(\uart/uart_idr_t [6]),
    .i12(\uart/uart_idr_t [6]),
    .i13(\uart/uart_idr_t [6]),
    .i14(\uart/uart_idr_t [6]),
    .i15(\uart/uart_idr_t [6]),
    .i2(\uart/n78 [6]),
    .i3(\uart/n78 [6]),
    .i4(\uart/n78 [6]),
    .i5(\uart/n78 [6]),
    .i6(\uart/n78 [6]),
    .i7(\uart/n78 [6]),
    .i8(\uart/n78 [6]),
    .i9(\uart/n78 [6]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n106 [6]));  // ../src/uart.v(261)
  binary_mux_s4_w1 \uart/mux47_b7  (
    .i0(\uart/n45 [7]),
    .i1(\uart/uart_idr_t [7]),
    .i10(\uart/uart_idr_t [7]),
    .i11(\uart/uart_idr_t [7]),
    .i12(\uart/uart_idr_t [7]),
    .i13(\uart/uart_idr_t [7]),
    .i14(\uart/uart_idr_t [7]),
    .i15(\uart/uart_idr_t [7]),
    .i2(\uart/n78 [7]),
    .i3(\uart/n78 [7]),
    .i4(\uart/n78 [7]),
    .i5(\uart/n78 [7]),
    .i6(\uart/n78 [7]),
    .i7(\uart/n78 [7]),
    .i8(\uart/n78 [7]),
    .i9(\uart/n78 [7]),
    .sel(\uart/uart_status_rxd ),
    .o(\uart/n106 [7]));  // ../src/uart.v(261)
  and \uart/mux4_sel_is_3  (\uart/mux4_sel_is_3_o , mem_la_addr[2], mem_la_addr[3]);
  and \uart/mux51_b0_sel_is_3  (\uart/mux51_b0_sel_is_3_o , \uart/uart_op_clock , \uart/mux44_b0_sel_is_26_o );
  binary_mux_s1_w1 \uart/mux53_b0  (
    .i0(\uart/uart_status_txd [0]),
    .i1(1'b1),
    .sel(\uart/uart_op_clock_by_3 ),
    .o(\uart/n31 [0]));  // ../src/uart.v(139)
  binary_mux_s1_w1 \uart/mux53_b1  (
    .i0(\uart/uart_status_txd [1]),
    .i1(1'b0),
    .sel(\uart/uart_op_clock_by_3 ),
    .o(\uart/n31 [1]));  // ../src/uart.v(139)
  binary_mux_s1_w1 \uart/mux53_b10  (
    .i0(\uart/uart_status_txd [2]),
    .i1(\uart/n35 [2]),
    .sel(\uart/uart_op_clock_by_3 ),
    .o(\uart/n36 [2]));  // ../src/uart.v(139)
  binary_mux_s1_w1 \uart/mux53_b11  (
    .i0(\uart/uart_status_txd [3]),
    .i1(\uart/n35 [3]),
    .sel(\uart/uart_op_clock_by_3 ),
    .o(\uart/n36 [3]));  // ../src/uart.v(139)
  binary_mux_s1_w1 \uart/mux53_b12  (
    .i0(\uart/uart_status_txd [0]),
    .i1(1'b0),
    .sel(\uart/uart_op_clock_by_3 ),
    .o(\uart/n37 [0]));  // ../src/uart.v(139)
  binary_mux_s1_w1 \uart/mux53_b14  (
    .i0(\uart/uart_status_txd [2]),
    .i1(1'b0),
    .sel(\uart/uart_op_clock_by_3 ),
    .o(\uart/n37 [2]));  // ../src/uart.v(139)
  binary_mux_s1_w1 \uart/mux53_b15  (
    .i0(\uart/uart_status_txd [3]),
    .i1(1'b0),
    .sel(\uart/uart_op_clock_by_3 ),
    .o(\uart/n37 [3]));  // ../src/uart.v(139)
  binary_mux_s1_w1 \uart/mux53_b5  (
    .i0(\uart/uart_status_txd [1]),
    .i1(1'b1),
    .sel(\uart/uart_op_clock_by_3 ),
    .o(\uart/n32 [1]));  // ../src/uart.v(139)
  binary_mux_s1_w1 \uart/mux53_b8  (
    .i0(\uart/uart_status_txd [0]),
    .i1(\uart/n35 [0]),
    .sel(\uart/uart_op_clock_by_3 ),
    .o(\uart/n36 [0]));  // ../src/uart.v(139)
  binary_mux_s1_w1 \uart/mux53_b9  (
    .i0(\uart/uart_status_txd [1]),
    .i1(\uart/n35 [1]),
    .sel(\uart/uart_op_clock_by_3 ),
    .o(\uart/n36 [1]));  // ../src/uart.v(139)
  and \uart/mux5_b0_sel_is_2  (\uart/mux5_b0_sel_is_2_o , mem_la_addr$2$_neg, mem_la_addr[3]);
  and \uart/mux6_b0_sel_is_4  (\uart/mux6_b0_sel_is_4_o , mem_la_addr$2$_neg, mem_la_addr$3$_neg, \uart/n9 );
  binary_mux_s2_w1 \uart/mux8_b0  (
    .i0(\uart/uart_odr [0]),
    .i1(\uart/uart_idr [0]),
    .i2(\uart/uart_bsrr [0]),
    .i3(\uart/uart_sr [0]),
    .sel(mem_la_addr[3:2]),
    .o(\uart/n16 [0]));  // ../src/uart.v(100)
  binary_mux_s2_w1 \uart/mux8_b1  (
    .i0(\uart/uart_odr [1]),
    .i1(\uart/uart_idr [1]),
    .i2(\uart/uart_bsrr [1]),
    .i3(\uart/uart_status_rx ),
    .sel(mem_la_addr[3:2]),
    .o(\uart/n16 [1]));  // ../src/uart.v(100)
  AL_MUX \uart/mux8_b10  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [10]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [10]));
  AL_MUX \uart/mux8_b11  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [11]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [11]));
  AL_MUX \uart/mux8_b12  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [12]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [12]));
  AL_MUX \uart/mux8_b13  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [13]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [13]));
  AL_MUX \uart/mux8_b14  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [14]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [14]));
  AL_MUX \uart/mux8_b15  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [15]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [15]));
  AL_MUX \uart/mux8_b16  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [16]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [16]));
  AL_MUX \uart/mux8_b17  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [17]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [17]));
  AL_MUX \uart/mux8_b18  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [18]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [18]));
  AL_MUX \uart/mux8_b19  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [19]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [19]));
  binary_mux_s2_w1 \uart/mux8_b2  (
    .i0(\uart/uart_odr [2]),
    .i1(\uart/uart_idr [2]),
    .i2(\uart/uart_bsrr [2]),
    .i3(\uart/uart_status_fe ),
    .sel(mem_la_addr[3:2]),
    .o(\uart/n16 [2]));  // ../src/uart.v(100)
  AL_MUX \uart/mux8_b20  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [20]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [20]));
  AL_MUX \uart/mux8_b21  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [21]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [21]));
  AL_MUX \uart/mux8_b22  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [22]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [22]));
  AL_MUX \uart/mux8_b23  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [23]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [23]));
  AL_MUX \uart/mux8_b24  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [24]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [24]));
  AL_MUX \uart/mux8_b25  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [25]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [25]));
  AL_MUX \uart/mux8_b26  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [26]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [26]));
  AL_MUX \uart/mux8_b27  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [27]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [27]));
  AL_MUX \uart/mux8_b28  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [28]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [28]));
  AL_MUX \uart/mux8_b29  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [29]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [29]));
  binary_mux_s2_w1 \uart/mux8_b3  (
    .i0(\uart/uart_odr [3]),
    .i1(\uart/uart_idr [3]),
    .i2(\uart/uart_bsrr [3]),
    .i3(1'b0),
    .sel(mem_la_addr[3:2]),
    .o(\uart/n16 [3]));  // ../src/uart.v(100)
  AL_MUX \uart/mux8_b30  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [30]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [30]));
  AL_MUX \uart/mux8_b31  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [31]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [31]));
  binary_mux_s2_w1 \uart/mux8_b4  (
    .i0(\uart/uart_odr [4]),
    .i1(\uart/uart_idr [4]),
    .i2(\uart/uart_bsrr [4]),
    .i3(1'b0),
    .sel(mem_la_addr[3:2]),
    .o(\uart/n16 [4]));  // ../src/uart.v(100)
  binary_mux_s2_w1 \uart/mux8_b5  (
    .i0(\uart/uart_odr [5]),
    .i1(\uart/uart_idr [5]),
    .i2(\uart/uart_bsrr [5]),
    .i3(1'b0),
    .sel(mem_la_addr[3:2]),
    .o(\uart/n16 [5]));  // ../src/uart.v(100)
  binary_mux_s2_w1 \uart/mux8_b6  (
    .i0(\uart/uart_odr [6]),
    .i1(\uart/uart_idr [6]),
    .i2(\uart/uart_bsrr [6]),
    .i3(1'b0),
    .sel(mem_la_addr[3:2]),
    .o(\uart/n16 [6]));  // ../src/uart.v(100)
  binary_mux_s2_w1 \uart/mux8_b7  (
    .i0(\uart/uart_odr [7]),
    .i1(\uart/uart_idr [7]),
    .i2(\uart/uart_bsrr [7]),
    .i3(1'b0),
    .sel(mem_la_addr[3:2]),
    .o(\uart/n16 [7]));  // ../src/uart.v(100)
  AL_MUX \uart/mux8_b8  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [8]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [8]));
  AL_MUX \uart/mux8_b9  (
    .i0(1'b0),
    .i1(\uart/uart_bsrr [9]),
    .sel(\uart/mux5_b0_sel_is_2_o ),
    .o(\uart/n16 [9]));
  and \uart/mux9_b0_sel_is_3  (\uart/mux9_b0_sel_is_3_o , mem_la_write, \uart/mux5_b0_sel_is_2_o );
  ne_w4 \uart/neq0  (
    .i0(\uart/uart_status_txd ),
    .i1(4'b0000),
    .o(\uart/n0 ));  // ../src/uart.v(42)
  reg_ar_as_w1 \uart/reg0_b0  (
    .clk(clk),
    .d(\uart/n16 [0]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[0]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b1  (
    .clk(clk),
    .d(\uart/n16 [1]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[1]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b10  (
    .clk(clk),
    .d(\uart/n16 [10]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[10]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b11  (
    .clk(clk),
    .d(\uart/n16 [11]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[11]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b12  (
    .clk(clk),
    .d(\uart/n16 [12]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[12]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b13  (
    .clk(clk),
    .d(\uart/n16 [13]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[13]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b14  (
    .clk(clk),
    .d(\uart/n16 [14]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[14]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b15  (
    .clk(clk),
    .d(\uart/n16 [15]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[15]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b16  (
    .clk(clk),
    .d(\uart/n16 [16]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[16]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b17  (
    .clk(clk),
    .d(\uart/n16 [17]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[17]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b18  (
    .clk(clk),
    .d(\uart/n16 [18]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[18]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b19  (
    .clk(clk),
    .d(\uart/n16 [19]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[19]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b2  (
    .clk(clk),
    .d(\uart/n16 [2]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[2]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b20  (
    .clk(clk),
    .d(\uart/n16 [20]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[20]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b21  (
    .clk(clk),
    .d(\uart/n16 [21]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[21]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b22  (
    .clk(clk),
    .d(\uart/n16 [22]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[22]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b23  (
    .clk(clk),
    .d(\uart/n16 [23]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[23]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b24  (
    .clk(clk),
    .d(\uart/n16 [24]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[24]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b25  (
    .clk(clk),
    .d(\uart/n16 [25]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[25]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b26  (
    .clk(clk),
    .d(\uart/n16 [26]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[26]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b27  (
    .clk(clk),
    .d(\uart/n16 [27]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[27]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b28  (
    .clk(clk),
    .d(\uart/n16 [28]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[28]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b29  (
    .clk(clk),
    .d(\uart/n16 [29]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[29]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b3  (
    .clk(clk),
    .d(\uart/n16 [3]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[3]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b30  (
    .clk(clk),
    .d(\uart/n16 [30]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[30]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b31  (
    .clk(clk),
    .d(\uart/n16 [31]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[31]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b4  (
    .clk(clk),
    .d(\uart/n16 [4]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[4]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b5  (
    .clk(clk),
    .d(\uart/n16 [5]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[5]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b6  (
    .clk(clk),
    .d(\uart/n16 [6]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[6]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b7  (
    .clk(clk),
    .d(\uart/n16 [7]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[7]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b8  (
    .clk(clk),
    .d(\uart/n16 [8]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[8]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg0_b9  (
    .clk(clk),
    .d(\uart/n16 [9]),
    .en(\uart/mux14_b0_sel_is_1_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(uart_do[9]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg10_b0  (
    .clk(clk),
    .d(\uart/n4 [0]),
    .en(\uart/n2 ),
    .reset(1'b0),
    .set(~resetn),
    .q(\uart/uart_op_clock_by_3_c [0]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg10_b1  (
    .clk(clk),
    .d(\uart/n4 [1]),
    .en(\uart/n2 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_op_clock_by_3_c [1]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b0  (
    .clk(clk),
    .d(\uart/n6 [0]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [0]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b1  (
    .clk(clk),
    .d(\uart/n6 [1]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [1]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b10  (
    .clk(clk),
    .d(\uart/n6 [10]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [10]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b11  (
    .clk(clk),
    .d(\uart/n6 [11]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [11]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b12  (
    .clk(clk),
    .d(\uart/n6 [12]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [12]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b13  (
    .clk(clk),
    .d(\uart/n6 [13]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [13]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b14  (
    .clk(clk),
    .d(\uart/n6 [14]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [14]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b15  (
    .clk(clk),
    .d(\uart/n6 [15]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [15]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b16  (
    .clk(clk),
    .d(\uart/n6 [16]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [16]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b17  (
    .clk(clk),
    .d(\uart/n6 [17]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [17]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b18  (
    .clk(clk),
    .d(\uart/n6 [18]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [18]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b19  (
    .clk(clk),
    .d(\uart/n6 [19]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [19]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b2  (
    .clk(clk),
    .d(\uart/n6 [2]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [2]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b20  (
    .clk(clk),
    .d(\uart/n6 [20]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [20]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b21  (
    .clk(clk),
    .d(\uart/n6 [21]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [21]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b22  (
    .clk(clk),
    .d(\uart/n6 [22]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [22]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b23  (
    .clk(clk),
    .d(\uart/n6 [23]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [23]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b24  (
    .clk(clk),
    .d(\uart/n6 [24]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [24]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b25  (
    .clk(clk),
    .d(\uart/n6 [25]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [25]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b26  (
    .clk(clk),
    .d(\uart/n6 [26]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [26]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b27  (
    .clk(clk),
    .d(\uart/n6 [27]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [27]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b28  (
    .clk(clk),
    .d(\uart/n6 [28]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [28]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b29  (
    .clk(clk),
    .d(\uart/n6 [29]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [29]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b3  (
    .clk(clk),
    .d(\uart/n6 [3]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [3]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b30  (
    .clk(clk),
    .d(\uart/n6 [30]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [30]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b31  (
    .clk(clk),
    .d(\uart/n6 [31]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [31]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b4  (
    .clk(clk),
    .d(\uart/n6 [4]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [4]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b5  (
    .clk(clk),
    .d(\uart/n6 [5]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [5]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b6  (
    .clk(clk),
    .d(\uart/n6 [6]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [6]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b7  (
    .clk(clk),
    .d(\uart/n6 [7]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [7]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b8  (
    .clk(clk),
    .d(\uart/n6 [8]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [8]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg1_b9  (
    .clk(clk),
    .d(\uart/n6 [9]),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_counter [9]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b0  (
    .clk(clk),
    .d(mem_la_wdata[0]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [0]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b1  (
    .clk(clk),
    .d(mem_la_wdata[1]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(~resetn),
    .q(\uart/uart_bsrr [1]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b10  (
    .clk(clk),
    .d(mem_la_wdata[10]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [10]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b11  (
    .clk(clk),
    .d(mem_la_wdata[11]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [11]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b12  (
    .clk(clk),
    .d(mem_la_wdata[12]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [12]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b13  (
    .clk(clk),
    .d(mem_la_wdata[13]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [13]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b14  (
    .clk(clk),
    .d(mem_la_wdata[14]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [14]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b15  (
    .clk(clk),
    .d(mem_la_wdata[15]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [15]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b16  (
    .clk(clk),
    .d(mem_la_wdata[16]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [16]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b17  (
    .clk(clk),
    .d(mem_la_wdata[17]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [17]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b18  (
    .clk(clk),
    .d(mem_la_wdata[18]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [18]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b19  (
    .clk(clk),
    .d(mem_la_wdata[19]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [19]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b2  (
    .clk(clk),
    .d(mem_la_wdata[2]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [2]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b20  (
    .clk(clk),
    .d(mem_la_wdata[20]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [20]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b21  (
    .clk(clk),
    .d(mem_la_wdata[21]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [21]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b22  (
    .clk(clk),
    .d(mem_la_wdata[22]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [22]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b23  (
    .clk(clk),
    .d(mem_la_wdata[23]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [23]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b24  (
    .clk(clk),
    .d(mem_la_wdata[24]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [24]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b25  (
    .clk(clk),
    .d(mem_la_wdata[25]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [25]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b26  (
    .clk(clk),
    .d(mem_la_wdata[26]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [26]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b27  (
    .clk(clk),
    .d(mem_la_wdata[27]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [27]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b28  (
    .clk(clk),
    .d(mem_la_wdata[28]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [28]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b29  (
    .clk(clk),
    .d(mem_la_wdata[29]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [29]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b3  (
    .clk(clk),
    .d(mem_la_wdata[3]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [3]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b30  (
    .clk(clk),
    .d(mem_la_wdata[30]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [30]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b31  (
    .clk(clk),
    .d(mem_la_wdata[31]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [31]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b4  (
    .clk(clk),
    .d(mem_la_wdata[4]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [4]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b5  (
    .clk(clk),
    .d(mem_la_wdata[5]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [5]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b6  (
    .clk(clk),
    .d(mem_la_wdata[6]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [6]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b7  (
    .clk(clk),
    .d(mem_la_wdata[7]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [7]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b8  (
    .clk(clk),
    .d(mem_la_wdata[8]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [8]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg2_b9  (
    .clk(clk),
    .d(mem_la_wdata[9]),
    .en(\uart/mux12_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_bsrr [9]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg3_b0  (
    .clk(clk),
    .d(mem_la_wdata[0]),
    .en(\uart/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\uart/uart_odr [0]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg3_b1  (
    .clk(clk),
    .d(mem_la_wdata[1]),
    .en(\uart/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\uart/uart_odr [1]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg3_b2  (
    .clk(clk),
    .d(mem_la_wdata[2]),
    .en(\uart/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\uart/uart_odr [2]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg3_b3  (
    .clk(clk),
    .d(mem_la_wdata[3]),
    .en(\uart/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\uart/uart_odr [3]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg3_b4  (
    .clk(clk),
    .d(mem_la_wdata[4]),
    .en(\uart/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\uart/uart_odr [4]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg3_b5  (
    .clk(clk),
    .d(mem_la_wdata[5]),
    .en(\uart/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\uart/uart_odr [5]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg3_b6  (
    .clk(clk),
    .d(mem_la_wdata[6]),
    .en(\uart/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\uart/uart_odr [6]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg3_b7  (
    .clk(clk),
    .d(mem_la_wdata[7]),
    .en(\uart/mux15_b0_sel_is_2_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\uart/uart_odr [7]));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/reg4_b0  (
    .clk(clk),
    .d(\uart/n38 [0]),
    .en(\uart/n30 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_status_txd [0]));  // ../src/uart.v(145)
  reg_ar_as_w1 \uart/reg4_b1  (
    .clk(clk),
    .d(\uart/n38 [1]),
    .en(\uart/n30 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_status_txd [1]));  // ../src/uart.v(145)
  reg_ar_as_w1 \uart/reg4_b2  (
    .clk(clk),
    .d(\uart/n38 [2]),
    .en(\uart/n30 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_status_txd [2]));  // ../src/uart.v(145)
  reg_ar_as_w1 \uart/reg4_b3  (
    .clk(clk),
    .d(\uart/n38 [3]),
    .en(\uart/n30 ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_status_txd [3]));  // ../src/uart.v(145)
  reg_ar_as_w1 \uart/reg5_b0  (
    .clk(clk),
    .d(\uart/n100 [0]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_status_rxd [0]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg5_b1  (
    .clk(clk),
    .d(\uart/n100 [1]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_status_rxd [1]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg5_b2  (
    .clk(clk),
    .d(\uart/n100 [2]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_status_rxd [2]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg5_b3  (
    .clk(clk),
    .d(\uart/n100 [3]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_status_rxd [3]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg6_b0  (
    .clk(clk),
    .d(\uart/uart_idr_t [0]),
    .en(\uart/mux51_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr [0]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg6_b1  (
    .clk(clk),
    .d(\uart/uart_idr_t [1]),
    .en(\uart/mux51_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr [1]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg6_b2  (
    .clk(clk),
    .d(\uart/uart_idr_t [2]),
    .en(\uart/mux51_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr [2]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg6_b3  (
    .clk(clk),
    .d(\uart/uart_idr_t [3]),
    .en(\uart/mux51_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr [3]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg6_b4  (
    .clk(clk),
    .d(\uart/uart_idr_t [4]),
    .en(\uart/mux51_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr [4]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg6_b5  (
    .clk(clk),
    .d(\uart/uart_idr_t [5]),
    .en(\uart/mux51_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr [5]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg6_b6  (
    .clk(clk),
    .d(\uart/uart_idr_t [6]),
    .en(\uart/mux51_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr [6]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg6_b7  (
    .clk(clk),
    .d(\uart/uart_idr_t [7]),
    .en(\uart/mux51_b0_sel_is_3_o ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr [7]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg7_b0  (
    .clk(clk),
    .d(\uart/n106 [0]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr_t [0]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg7_b1  (
    .clk(clk),
    .d(\uart/n106 [1]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr_t [1]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg7_b2  (
    .clk(clk),
    .d(\uart/n106 [2]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr_t [2]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg7_b3  (
    .clk(clk),
    .d(\uart/n106 [3]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr_t [3]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg7_b4  (
    .clk(clk),
    .d(\uart/n106 [4]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr_t [4]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg7_b5  (
    .clk(clk),
    .d(\uart/n106 [5]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr_t [5]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg7_b6  (
    .clk(clk),
    .d(\uart/n106 [6]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr_t [6]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg7_b7  (
    .clk(clk),
    .d(\uart/n106 [7]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_idr_t [7]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg8_b0  (
    .clk(clk),
    .d(\uart/n102 [0]),
    .en(\uart/uart_op_clock ),
    .reset(1'b0),
    .set(~resetn),
    .q(\uart/uart_cnt_rx [0]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg8_b1  (
    .clk(clk),
    .d(\uart/n102 [1]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_cnt_rx [1]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg8_b2  (
    .clk(clk),
    .d(\uart/n102 [2]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_cnt_rx [2]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg9_b0  (
    .clk(clk),
    .d(\uart/n101 [0]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_smp_rx [0]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg9_b1  (
    .clk(clk),
    .d(\uart/n101 [1]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_smp_rx [1]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg9_b2  (
    .clk(clk),
    .d(\uart/n101 [2]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_smp_rx [2]));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/reg9_b3  (
    .clk(clk),
    .d(\uart/n101 [3]),
    .en(\uart/uart_op_clock ),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_smp_rx [3]));  // ../src/uart.v(263)
  add_pu3_mu3_o3 \uart/sub0  (
    .i0(\uart/uart_status_txd [2:0]),
    .i1(3'b010),
    .o(\uart/n33 [2:0]));  // ../src/uart.v(131)
  add_pu4_mu4_o5 \uart/sub1  (
    .i0(\uart/uart_status_rxd ),
    .i1(4'b0010),
    .o(\uart/n57 ));  // ../src/uart.v(222)
  reg_ar_as_w1 \uart/txd_o_reg  (
    .clk(clk),
    .d(\uart/n39 ),
    .en(\uart/n30 ),
    .reset(1'b0),
    .set(~resetn),
    .q(txd));  // ../src/uart.v(145)
  or \uart/u12  (\uart/n3 , \uart/uart_op_clock_by_3_c [0], \uart/uart_op_clock_by_3_c [1]);  // ../src/uart.v(63)
  or \uart/u13  (\uart/n30 , \uart/n29 , \uart/uart_trigger_tx );  // ../src/uart.v(114)
  or \uart/u14  (\uart/n83 , \uart/uart_status_txd [0], \uart/uart_status_txd [1]);  // ../src/uart.v(114)
  AL_MUX \uart/u17  (
    .i0(\uart/uart_status_fe ),
    .i1(1'b0),
    .sel(\uart/uart_status_rx_clr ),
    .o(\uart/n43 ));  // ../src/uart.v(176)
  not \uart/u18  (\uart/n44 , rxd);  // ../src/uart.v(182)
  and \uart/u19  (\uart/n59 [0], \uart/n87 , \uart/n96 );  // ../src/uart.v(222)
  and \uart/u2  (\uart/uart_op_clock_by_3 , \uart/uart_op_clock_by_3_c [0], \uart/uart_op_clock );  // ../src/uart.v(37)
  and \uart/u20  (\uart/n59 [4], \uart/n87 , \uart/n57 [2]);  // ../src/uart.v(222)
  or \uart/u22  (\uart/n56 , \uart/uart_cnt_rx [0], \uart/uart_cnt_rx [1]);  // ../src/uart.v(209)
  or \uart/u23  (\uart/n84 , \uart/n57 [3], \uart/n57 [4]);  // ../src/uart.v(222)
  and \uart/u24  (\uart/n60 , \uart/n59 [7], \uart/n58 );  // ../src/uart.v(222)
  and \uart/u25  (\uart/n85 , \uart/n57 [0], \uart/n97 );  // ../src/uart.v(222)
  and \uart/u26  (\uart/n62 , \uart/n59 [6], \uart/n58 );  // ../src/uart.v(222)
  and \uart/u27  (\uart/n86 , \uart/n57 [0], \uart/n57 [1]);  // ../src/uart.v(222)
  and \uart/u28  (\uart/n64 , \uart/n59 [5], \uart/n58 );  // ../src/uart.v(222)
  and \uart/u29  (\uart/n87 , \uart/n89 , \uart/n97 );  // ../src/uart.v(222)
  or \uart/u3  (\uart/uart_sr [0], \uart/n0 , \uart/uart_trigger_tx );  // ../src/uart.v(42)
  and \uart/u30  (\uart/n66 , \uart/n59 [4], \uart/n58 );  // ../src/uart.v(222)
  and \uart/u31  (\uart/n88 , \uart/n89 , \uart/n57 [1]);  // ../src/uart.v(222)
  and \uart/u32  (\uart/n68 , \uart/n59 [3], \uart/n58 );  // ../src/uart.v(222)
  not \uart/u33  (\uart/n96 , \uart/n57 [2]);  // ../src/uart.v(222)
  and \uart/u34  (\uart/n70 , \uart/n59 [2], \uart/n58 );  // ../src/uart.v(222)
  not \uart/u35  (\uart/n97 , \uart/n57 [1]);  // ../src/uart.v(222)
  and \uart/u36  (\uart/n72 , \uart/n59 [1], \uart/n58 );  // ../src/uart.v(222)
  or \uart/u37  (\uart/n91 , \uart/n99 , \uart/n98 );  // ../src/uart.v(250)
  and \uart/u38  (\uart/n74 , \uart/n59 [0], \uart/n58 );  // ../src/uart.v(222)
  or \uart/u39  (\uart/n98 , \uart/uart_smp_rx [2], \uart/uart_smp_rx [3]);  // ../src/uart.v(250)
  or \uart/u40  (\uart/n29 , \uart/n83 , \uart/n82 );  // ../src/uart.v(114)
  or \uart/u41  (\uart/n82 , \uart/uart_status_txd [2], \uart/uart_status_txd [3]);  // ../src/uart.v(114)
  not \uart/u48  (\uart/n58 , \uart/n84 );  // ../src/uart.v(222)
  or \uart/u49  (\uart/n99 , \uart/uart_smp_rx [0], \uart/uart_smp_rx [1]);  // ../src/uart.v(250)
  and \uart/u50  (\uart/n59 [3], \uart/n86 , \uart/n96 );  // ../src/uart.v(222)
  and \uart/u51  (\uart/n59 [7], \uart/n86 , \uart/n57 [2]);  // ../src/uart.v(222)
  and \uart/u52  (\uart/n59 [2], \uart/n88 , \uart/n96 );  // ../src/uart.v(222)
  and \uart/u53  (\uart/n59 [6], \uart/n88 , \uart/n57 [2]);  // ../src/uart.v(222)
  and \uart/u54  (\uart/n59 [1], \uart/n85 , \uart/n96 );  // ../src/uart.v(222)
  not \uart/u55  (\uart/n89 , \uart/n57 [0]);  // ../src/uart.v(222)
  and \uart/u58  (\uart/n59 [5], \uart/n85 , \uart/n57 [2]);  // ../src/uart.v(222)
  AL_MUX \uart/u60  (
    .i0(\uart/n43 ),
    .i1(\uart/n91 ),
    .sel(\uart/mux51_b0_sel_is_3_o ),
    .o(\uart/n112 ));
  and \uart/u7_sel_is_3  (\uart/u7_sel_is_3_o , mem_la_write, \uart/mux4_sel_is_3_o );
  and \uart/u9_sel_is_3  (\uart/u9_sel_is_3_o , uart_sel, \uart/u7_sel_is_3_o );
  reg_ar_as_w1 \uart/uart_op_clock_reg  (
    .clk(clk),
    .d(\uart/n2 ),
    .en(~\picorv32_core/n407 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\uart/uart_op_clock ));  // ../src/uart.v(102)
  reg_ar_as_w1 \uart/uart_status_fe_reg  (
    .clk(clk),
    .d(\uart/n112 ),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_status_fe ));  // ../src/uart.v(263)
  reg_ar_as_w1 \uart/uart_status_rx_clr_reg  (
    .clk(clk),
    .d(\uart/u9_sel_is_3_o ),
    .en(1'b1),
    .reset(~resetn),
    .set(1'b0),
    .q(\uart/uart_status_rx_clr ));  // ../src/uart.v(102)
  reg_ar_ss_w1 \uart/uart_status_rx_reg  (
    .clk(clk),
    .d(1'b0),
    .en(\uart/uart_status_rx_clr ),
    .reset(~resetn),
    .set(\uart/mux51_b0_sel_is_3_o ),
    .q(\uart/uart_status_rx ));  // ../src/uart.v(263)
  not \uart/uart_status_rxd[0]_inv  (\uart/uart_status_rxd$0$_neg , \uart/uart_status_rxd [0]);
  not \uart/uart_status_rxd[2]_inv  (\uart/uart_status_rxd$2$_neg , \uart/uart_status_rxd [2]);
  reg_ar_ss_w1 \uart/uart_trigger_tx_reg  (
    .clk(clk),
    .d(1'b0),
    .en(\uart/uart_op_clock_by_3 ),
    .reset(~resetn),
    .set(\uart/mux13_b0_sel_is_3_o ),
    .q(\uart/uart_trigger_tx ));  // ../src/uart.v(102)

endmodule 

module add_pu2_pu2_o2
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output [1:0] o;

  wire net_a0;
  wire net_a1;
  wire net_b0;
  wire net_b1;
  wire net_cout0;
  wire net_cout1;
  wire net_sum0;
  wire net_sum1;

  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));

endmodule 

module eq_w2
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output o;

  wire or_xor_i0$0$_i1$0$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;

  not none_diff (o, or_xor_i0$0$_i1$0$_o_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, xor_i0$1$_i1$1$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);

endmodule 

module eq_w20
  (
  i0,
  i1,
  o
  );

  input [19:0] i0;
  input [19:0] i1;
  output o;

  wire or_or_or_or_xor_i0$0_o;
  wire or_or_or_xor_i0$0$_i_o;
  wire or_or_or_xor_i0$10$__o;
  wire or_or_xor_i0$0$_i1$0_o;
  wire or_or_xor_i0$10$_i1$_o;
  wire or_or_xor_i0$15$_i1$_o;
  wire or_or_xor_i0$5$_i1$5_o;
  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$10$_i1$10$_o;
  wire or_xor_i0$12$_i1$12$_o;
  wire or_xor_i0$13$_i1$13$_o;
  wire or_xor_i0$15$_i1$15$_o;
  wire or_xor_i0$17$_i1$17$_o;
  wire or_xor_i0$18$_i1$18$_o;
  wire or_xor_i0$2$_i1$2$_o_o;
  wire or_xor_i0$3$_i1$3$_o_o;
  wire or_xor_i0$5$_i1$5$_o_o;
  wire or_xor_i0$7$_i1$7$_o_o;
  wire or_xor_i0$8$_i1$8$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$10$_i1$10$_o;
  wire xor_i0$11$_i1$11$_o;
  wire xor_i0$12$_i1$12$_o;
  wire xor_i0$13$_i1$13$_o;
  wire xor_i0$14$_i1$14$_o;
  wire xor_i0$15$_i1$15$_o;
  wire xor_i0$16$_i1$16$_o;
  wire xor_i0$17$_i1$17$_o;
  wire xor_i0$18$_i1$18$_o;
  wire xor_i0$19$_i1$19$_o;
  wire xor_i0$2$_i1$2$_o;
  wire xor_i0$3$_i1$3$_o;
  wire xor_i0$4$_i1$4$_o;
  wire xor_i0$5$_i1$5$_o;
  wire xor_i0$6$_i1$6$_o;
  wire xor_i0$7$_i1$7$_o;
  wire xor_i0$8$_i1$8$_o;
  wire xor_i0$9$_i1$9$_o;

  not none_diff (o, or_or_or_or_xor_i0$0_o);
  or or_or_or_or_xor_i0$0 (or_or_or_or_xor_i0$0_o, or_or_or_xor_i0$0$_i_o, or_or_or_xor_i0$10$__o);
  or or_or_or_xor_i0$0$_i (or_or_or_xor_i0$0$_i_o, or_or_xor_i0$0$_i1$0_o, or_or_xor_i0$5$_i1$5_o);
  or or_or_or_xor_i0$10$_ (or_or_or_xor_i0$10$__o, or_or_xor_i0$10$_i1$_o, or_or_xor_i0$15$_i1$_o);
  or or_or_xor_i0$0$_i1$0 (or_or_xor_i0$0$_i1$0_o, or_xor_i0$0$_i1$0$_o_o, or_xor_i0$2$_i1$2$_o_o);
  or or_or_xor_i0$10$_i1$ (or_or_xor_i0$10$_i1$_o, or_xor_i0$10$_i1$10$_o, or_xor_i0$12$_i1$12$_o);
  or or_or_xor_i0$15$_i1$ (or_or_xor_i0$15$_i1$_o, or_xor_i0$15$_i1$15$_o, or_xor_i0$17$_i1$17$_o);
  or or_or_xor_i0$5$_i1$5 (or_or_xor_i0$5$_i1$5_o, or_xor_i0$5$_i1$5$_o_o, or_xor_i0$7$_i1$7$_o_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, xor_i0$1$_i1$1$_o);
  or or_xor_i0$10$_i1$10$ (or_xor_i0$10$_i1$10$_o, xor_i0$10$_i1$10$_o, xor_i0$11$_i1$11$_o);
  or or_xor_i0$12$_i1$12$ (or_xor_i0$12$_i1$12$_o, xor_i0$12$_i1$12$_o, or_xor_i0$13$_i1$13$_o);
  or or_xor_i0$13$_i1$13$ (or_xor_i0$13$_i1$13$_o, xor_i0$13$_i1$13$_o, xor_i0$14$_i1$14$_o);
  or or_xor_i0$15$_i1$15$ (or_xor_i0$15$_i1$15$_o, xor_i0$15$_i1$15$_o, xor_i0$16$_i1$16$_o);
  or or_xor_i0$17$_i1$17$ (or_xor_i0$17$_i1$17$_o, xor_i0$17$_i1$17$_o, or_xor_i0$18$_i1$18$_o);
  or or_xor_i0$18$_i1$18$ (or_xor_i0$18$_i1$18$_o, xor_i0$18$_i1$18$_o, xor_i0$19$_i1$19$_o);
  or or_xor_i0$2$_i1$2$_o (or_xor_i0$2$_i1$2$_o_o, xor_i0$2$_i1$2$_o, or_xor_i0$3$_i1$3$_o_o);
  or or_xor_i0$3$_i1$3$_o (or_xor_i0$3$_i1$3$_o_o, xor_i0$3$_i1$3$_o, xor_i0$4$_i1$4$_o);
  or or_xor_i0$5$_i1$5$_o (or_xor_i0$5$_i1$5$_o_o, xor_i0$5$_i1$5$_o, xor_i0$6$_i1$6$_o);
  or or_xor_i0$7$_i1$7$_o (or_xor_i0$7$_i1$7$_o_o, xor_i0$7$_i1$7$_o, or_xor_i0$8$_i1$8$_o_o);
  or or_xor_i0$8$_i1$8$_o (or_xor_i0$8$_i1$8$_o_o, xor_i0$8$_i1$8$_o, xor_i0$9$_i1$9$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (xor_i0$10$_i1$10$_o, i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (xor_i0$11$_i1$11$_o, i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (xor_i0$12$_i1$12$_o, i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (xor_i0$13$_i1$13$_o, i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (xor_i0$14$_i1$14$_o, i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (xor_i0$15$_i1$15$_o, i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (xor_i0$16$_i1$16$_o, i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (xor_i0$17$_i1$17$_o, i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (xor_i0$18$_i1$18$_o, i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (xor_i0$19$_i1$19$_o, i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (xor_i0$3$_i1$3$_o, i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (xor_i0$4$_i1$4$_o, i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (xor_i0$5$_i1$5$_o, i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (xor_i0$6$_i1$6$_o, i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (xor_i0$7$_i1$7$_o, i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (xor_i0$8$_i1$8$_o, i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (xor_i0$9$_i1$9$_o, i0[9], i1[9]);

endmodule 

module eq_w28
  (
  i0,
  i1,
  o
  );

  input [27:0] i0;
  input [27:0] i1;
  output o;

  wire or_or_or_or_xor_i0$0_o;
  wire or_or_or_xor_i0$0$_i_o;
  wire or_or_or_xor_i0$14$__o;
  wire or_or_xor_i0$0$_i1$0_o;
  wire or_or_xor_i0$10$_i1$_o;
  wire or_or_xor_i0$14$_i1$_o;
  wire or_or_xor_i0$17$_i1$_o;
  wire or_or_xor_i0$21$_i1$_o;
  wire or_or_xor_i0$24$_i1$_o;
  wire or_or_xor_i0$3$_i1$3_o;
  wire or_or_xor_i0$7$_i1$7_o;
  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$1$_i1$1$_o_o;
  wire or_xor_i0$10$_i1$10$_o;
  wire or_xor_i0$12$_i1$12$_o;
  wire or_xor_i0$14$_i1$14$_o;
  wire or_xor_i0$15$_i1$15$_o;
  wire or_xor_i0$17$_i1$17$_o;
  wire or_xor_i0$19$_i1$19$_o;
  wire or_xor_i0$21$_i1$21$_o;
  wire or_xor_i0$22$_i1$22$_o;
  wire or_xor_i0$24$_i1$24$_o;
  wire or_xor_i0$26$_i1$26$_o;
  wire or_xor_i0$3$_i1$3$_o_o;
  wire or_xor_i0$5$_i1$5$_o_o;
  wire or_xor_i0$7$_i1$7$_o_o;
  wire or_xor_i0$8$_i1$8$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$10$_i1$10$_o;
  wire xor_i0$11$_i1$11$_o;
  wire xor_i0$12$_i1$12$_o;
  wire xor_i0$13$_i1$13$_o;
  wire xor_i0$14$_i1$14$_o;
  wire xor_i0$15$_i1$15$_o;
  wire xor_i0$16$_i1$16$_o;
  wire xor_i0$17$_i1$17$_o;
  wire xor_i0$18$_i1$18$_o;
  wire xor_i0$19$_i1$19$_o;
  wire xor_i0$2$_i1$2$_o;
  wire xor_i0$20$_i1$20$_o;
  wire xor_i0$21$_i1$21$_o;
  wire xor_i0$22$_i1$22$_o;
  wire xor_i0$23$_i1$23$_o;
  wire xor_i0$24$_i1$24$_o;
  wire xor_i0$25$_i1$25$_o;
  wire xor_i0$26$_i1$26$_o;
  wire xor_i0$27$_i1$27$_o;
  wire xor_i0$3$_i1$3$_o;
  wire xor_i0$4$_i1$4$_o;
  wire xor_i0$5$_i1$5$_o;
  wire xor_i0$6$_i1$6$_o;
  wire xor_i0$7$_i1$7$_o;
  wire xor_i0$8$_i1$8$_o;
  wire xor_i0$9$_i1$9$_o;

  not none_diff (o, or_or_or_or_xor_i0$0_o);
  or or_or_or_or_xor_i0$0 (or_or_or_or_xor_i0$0_o, or_or_or_xor_i0$0$_i_o, or_or_or_xor_i0$14$__o);
  or or_or_or_xor_i0$0$_i (or_or_or_xor_i0$0$_i_o, or_or_xor_i0$0$_i1$0_o, or_or_xor_i0$7$_i1$7_o);
  or or_or_or_xor_i0$14$_ (or_or_or_xor_i0$14$__o, or_or_xor_i0$14$_i1$_o, or_or_xor_i0$21$_i1$_o);
  or or_or_xor_i0$0$_i1$0 (or_or_xor_i0$0$_i1$0_o, or_xor_i0$0$_i1$0$_o_o, or_or_xor_i0$3$_i1$3_o);
  or or_or_xor_i0$10$_i1$ (or_or_xor_i0$10$_i1$_o, or_xor_i0$10$_i1$10$_o, or_xor_i0$12$_i1$12$_o);
  or or_or_xor_i0$14$_i1$ (or_or_xor_i0$14$_i1$_o, or_xor_i0$14$_i1$14$_o, or_or_xor_i0$17$_i1$_o);
  or or_or_xor_i0$17$_i1$ (or_or_xor_i0$17$_i1$_o, or_xor_i0$17$_i1$17$_o, or_xor_i0$19$_i1$19$_o);
  or or_or_xor_i0$21$_i1$ (or_or_xor_i0$21$_i1$_o, or_xor_i0$21$_i1$21$_o, or_or_xor_i0$24$_i1$_o);
  or or_or_xor_i0$24$_i1$ (or_or_xor_i0$24$_i1$_o, or_xor_i0$24$_i1$24$_o, or_xor_i0$26$_i1$26$_o);
  or or_or_xor_i0$3$_i1$3 (or_or_xor_i0$3$_i1$3_o, or_xor_i0$3$_i1$3$_o_o, or_xor_i0$5$_i1$5$_o_o);
  or or_or_xor_i0$7$_i1$7 (or_or_xor_i0$7$_i1$7_o, or_xor_i0$7$_i1$7$_o_o, or_or_xor_i0$10$_i1$_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, or_xor_i0$1$_i1$1$_o_o);
  or or_xor_i0$1$_i1$1$_o (or_xor_i0$1$_i1$1$_o_o, xor_i0$1$_i1$1$_o, xor_i0$2$_i1$2$_o);
  or or_xor_i0$10$_i1$10$ (or_xor_i0$10$_i1$10$_o, xor_i0$10$_i1$10$_o, xor_i0$11$_i1$11$_o);
  or or_xor_i0$12$_i1$12$ (or_xor_i0$12$_i1$12$_o, xor_i0$12$_i1$12$_o, xor_i0$13$_i1$13$_o);
  or or_xor_i0$14$_i1$14$ (or_xor_i0$14$_i1$14$_o, xor_i0$14$_i1$14$_o, or_xor_i0$15$_i1$15$_o);
  or or_xor_i0$15$_i1$15$ (or_xor_i0$15$_i1$15$_o, xor_i0$15$_i1$15$_o, xor_i0$16$_i1$16$_o);
  or or_xor_i0$17$_i1$17$ (or_xor_i0$17$_i1$17$_o, xor_i0$17$_i1$17$_o, xor_i0$18$_i1$18$_o);
  or or_xor_i0$19$_i1$19$ (or_xor_i0$19$_i1$19$_o, xor_i0$19$_i1$19$_o, xor_i0$20$_i1$20$_o);
  or or_xor_i0$21$_i1$21$ (or_xor_i0$21$_i1$21$_o, xor_i0$21$_i1$21$_o, or_xor_i0$22$_i1$22$_o);
  or or_xor_i0$22$_i1$22$ (or_xor_i0$22$_i1$22$_o, xor_i0$22$_i1$22$_o, xor_i0$23$_i1$23$_o);
  or or_xor_i0$24$_i1$24$ (or_xor_i0$24$_i1$24$_o, xor_i0$24$_i1$24$_o, xor_i0$25$_i1$25$_o);
  or or_xor_i0$26$_i1$26$ (or_xor_i0$26$_i1$26$_o, xor_i0$26$_i1$26$_o, xor_i0$27$_i1$27$_o);
  or or_xor_i0$3$_i1$3$_o (or_xor_i0$3$_i1$3$_o_o, xor_i0$3$_i1$3$_o, xor_i0$4$_i1$4$_o);
  or or_xor_i0$5$_i1$5$_o (or_xor_i0$5$_i1$5$_o_o, xor_i0$5$_i1$5$_o, xor_i0$6$_i1$6$_o);
  or or_xor_i0$7$_i1$7$_o (or_xor_i0$7$_i1$7$_o_o, xor_i0$7$_i1$7$_o, or_xor_i0$8$_i1$8$_o_o);
  or or_xor_i0$8$_i1$8$_o (or_xor_i0$8$_i1$8$_o_o, xor_i0$8$_i1$8$_o, xor_i0$9$_i1$9$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (xor_i0$10$_i1$10$_o, i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (xor_i0$11$_i1$11$_o, i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (xor_i0$12$_i1$12$_o, i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (xor_i0$13$_i1$13$_o, i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (xor_i0$14$_i1$14$_o, i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (xor_i0$15$_i1$15$_o, i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (xor_i0$16$_i1$16$_o, i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (xor_i0$17$_i1$17$_o, i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (xor_i0$18$_i1$18$_o, i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (xor_i0$19$_i1$19$_o, i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (xor_i0$20$_i1$20$_o, i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (xor_i0$21$_i1$21$_o, i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (xor_i0$22$_i1$22$_o, i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (xor_i0$23$_i1$23$_o, i0[23], i1[23]);
  xor \xor_i0[24]_i1[24]  (xor_i0$24$_i1$24$_o, i0[24], i1[24]);
  xor \xor_i0[25]_i1[25]  (xor_i0$25$_i1$25$_o, i0[25], i1[25]);
  xor \xor_i0[26]_i1[26]  (xor_i0$26$_i1$26$_o, i0[26], i1[26]);
  xor \xor_i0[27]_i1[27]  (xor_i0$27$_i1$27$_o, i0[27], i1[27]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (xor_i0$3$_i1$3$_o, i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (xor_i0$4$_i1$4$_o, i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (xor_i0$5$_i1$5$_o, i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (xor_i0$6$_i1$6$_o, i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (xor_i0$7$_i1$7$_o, i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (xor_i0$8$_i1$8$_o, i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (xor_i0$9$_i1$9$_o, i0[9], i1[9]);

endmodule 

module eq_w30
  (
  i0,
  i1,
  o
  );

  input [29:0] i0;
  input [29:0] i1;
  output o;

  wire or_or_or_or_xor_i0$0_o;
  wire or_or_or_xor_i0$0$_i_o;
  wire or_or_or_xor_i0$15$__o;
  wire or_or_or_xor_i0$22$__o;
  wire or_or_or_xor_i0$7$_i_o;
  wire or_or_xor_i0$0$_i1$0_o;
  wire or_or_xor_i0$11$_i1$_o;
  wire or_or_xor_i0$15$_i1$_o;
  wire or_or_xor_i0$18$_i1$_o;
  wire or_or_xor_i0$22$_i1$_o;
  wire or_or_xor_i0$26$_i1$_o;
  wire or_or_xor_i0$3$_i1$3_o;
  wire or_or_xor_i0$7$_i1$7_o;
  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$1$_i1$1$_o_o;
  wire or_xor_i0$11$_i1$11$_o;
  wire or_xor_i0$13$_i1$13$_o;
  wire or_xor_i0$15$_i1$15$_o;
  wire or_xor_i0$16$_i1$16$_o;
  wire or_xor_i0$18$_i1$18$_o;
  wire or_xor_i0$20$_i1$20$_o;
  wire or_xor_i0$22$_i1$22$_o;
  wire or_xor_i0$24$_i1$24$_o;
  wire or_xor_i0$26$_i1$26$_o;
  wire or_xor_i0$28$_i1$28$_o;
  wire or_xor_i0$3$_i1$3$_o_o;
  wire or_xor_i0$5$_i1$5$_o_o;
  wire or_xor_i0$7$_i1$7$_o_o;
  wire or_xor_i0$9$_i1$9$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$10$_i1$10$_o;
  wire xor_i0$11$_i1$11$_o;
  wire xor_i0$12$_i1$12$_o;
  wire xor_i0$13$_i1$13$_o;
  wire xor_i0$14$_i1$14$_o;
  wire xor_i0$15$_i1$15$_o;
  wire xor_i0$16$_i1$16$_o;
  wire xor_i0$17$_i1$17$_o;
  wire xor_i0$18$_i1$18$_o;
  wire xor_i0$19$_i1$19$_o;
  wire xor_i0$2$_i1$2$_o;
  wire xor_i0$20$_i1$20$_o;
  wire xor_i0$21$_i1$21$_o;
  wire xor_i0$22$_i1$22$_o;
  wire xor_i0$23$_i1$23$_o;
  wire xor_i0$24$_i1$24$_o;
  wire xor_i0$25$_i1$25$_o;
  wire xor_i0$26$_i1$26$_o;
  wire xor_i0$27$_i1$27$_o;
  wire xor_i0$28$_i1$28$_o;
  wire xor_i0$29$_i1$29$_o;
  wire xor_i0$3$_i1$3$_o;
  wire xor_i0$4$_i1$4$_o;
  wire xor_i0$5$_i1$5$_o;
  wire xor_i0$6$_i1$6$_o;
  wire xor_i0$7$_i1$7$_o;
  wire xor_i0$8$_i1$8$_o;
  wire xor_i0$9$_i1$9$_o;

  not none_diff (o, or_or_or_or_xor_i0$0_o);
  or or_or_or_or_xor_i0$0 (or_or_or_or_xor_i0$0_o, or_or_or_xor_i0$0$_i_o, or_or_or_xor_i0$15$__o);
  or or_or_or_xor_i0$0$_i (or_or_or_xor_i0$0$_i_o, or_or_xor_i0$0$_i1$0_o, or_or_or_xor_i0$7$_i_o);
  or or_or_or_xor_i0$15$_ (or_or_or_xor_i0$15$__o, or_or_xor_i0$15$_i1$_o, or_or_or_xor_i0$22$__o);
  or or_or_or_xor_i0$22$_ (or_or_or_xor_i0$22$__o, or_or_xor_i0$22$_i1$_o, or_or_xor_i0$26$_i1$_o);
  or or_or_or_xor_i0$7$_i (or_or_or_xor_i0$7$_i_o, or_or_xor_i0$7$_i1$7_o, or_or_xor_i0$11$_i1$_o);
  or or_or_xor_i0$0$_i1$0 (or_or_xor_i0$0$_i1$0_o, or_xor_i0$0$_i1$0$_o_o, or_or_xor_i0$3$_i1$3_o);
  or or_or_xor_i0$11$_i1$ (or_or_xor_i0$11$_i1$_o, or_xor_i0$11$_i1$11$_o, or_xor_i0$13$_i1$13$_o);
  or or_or_xor_i0$15$_i1$ (or_or_xor_i0$15$_i1$_o, or_xor_i0$15$_i1$15$_o, or_or_xor_i0$18$_i1$_o);
  or or_or_xor_i0$18$_i1$ (or_or_xor_i0$18$_i1$_o, or_xor_i0$18$_i1$18$_o, or_xor_i0$20$_i1$20$_o);
  or or_or_xor_i0$22$_i1$ (or_or_xor_i0$22$_i1$_o, or_xor_i0$22$_i1$22$_o, or_xor_i0$24$_i1$24$_o);
  or or_or_xor_i0$26$_i1$ (or_or_xor_i0$26$_i1$_o, or_xor_i0$26$_i1$26$_o, or_xor_i0$28$_i1$28$_o);
  or or_or_xor_i0$3$_i1$3 (or_or_xor_i0$3$_i1$3_o, or_xor_i0$3$_i1$3$_o_o, or_xor_i0$5$_i1$5$_o_o);
  or or_or_xor_i0$7$_i1$7 (or_or_xor_i0$7$_i1$7_o, or_xor_i0$7$_i1$7$_o_o, or_xor_i0$9$_i1$9$_o_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, or_xor_i0$1$_i1$1$_o_o);
  or or_xor_i0$1$_i1$1$_o (or_xor_i0$1$_i1$1$_o_o, xor_i0$1$_i1$1$_o, xor_i0$2$_i1$2$_o);
  or or_xor_i0$11$_i1$11$ (or_xor_i0$11$_i1$11$_o, xor_i0$11$_i1$11$_o, xor_i0$12$_i1$12$_o);
  or or_xor_i0$13$_i1$13$ (or_xor_i0$13$_i1$13$_o, xor_i0$13$_i1$13$_o, xor_i0$14$_i1$14$_o);
  or or_xor_i0$15$_i1$15$ (or_xor_i0$15$_i1$15$_o, xor_i0$15$_i1$15$_o, or_xor_i0$16$_i1$16$_o);
  or or_xor_i0$16$_i1$16$ (or_xor_i0$16$_i1$16$_o, xor_i0$16$_i1$16$_o, xor_i0$17$_i1$17$_o);
  or or_xor_i0$18$_i1$18$ (or_xor_i0$18$_i1$18$_o, xor_i0$18$_i1$18$_o, xor_i0$19$_i1$19$_o);
  or or_xor_i0$20$_i1$20$ (or_xor_i0$20$_i1$20$_o, xor_i0$20$_i1$20$_o, xor_i0$21$_i1$21$_o);
  or or_xor_i0$22$_i1$22$ (or_xor_i0$22$_i1$22$_o, xor_i0$22$_i1$22$_o, xor_i0$23$_i1$23$_o);
  or or_xor_i0$24$_i1$24$ (or_xor_i0$24$_i1$24$_o, xor_i0$24$_i1$24$_o, xor_i0$25$_i1$25$_o);
  or or_xor_i0$26$_i1$26$ (or_xor_i0$26$_i1$26$_o, xor_i0$26$_i1$26$_o, xor_i0$27$_i1$27$_o);
  or or_xor_i0$28$_i1$28$ (or_xor_i0$28$_i1$28$_o, xor_i0$28$_i1$28$_o, xor_i0$29$_i1$29$_o);
  or or_xor_i0$3$_i1$3$_o (or_xor_i0$3$_i1$3$_o_o, xor_i0$3$_i1$3$_o, xor_i0$4$_i1$4$_o);
  or or_xor_i0$5$_i1$5$_o (or_xor_i0$5$_i1$5$_o_o, xor_i0$5$_i1$5$_o, xor_i0$6$_i1$6$_o);
  or or_xor_i0$7$_i1$7$_o (or_xor_i0$7$_i1$7$_o_o, xor_i0$7$_i1$7$_o, xor_i0$8$_i1$8$_o);
  or or_xor_i0$9$_i1$9$_o (or_xor_i0$9$_i1$9$_o_o, xor_i0$9$_i1$9$_o, xor_i0$10$_i1$10$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (xor_i0$10$_i1$10$_o, i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (xor_i0$11$_i1$11$_o, i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (xor_i0$12$_i1$12$_o, i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (xor_i0$13$_i1$13$_o, i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (xor_i0$14$_i1$14$_o, i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (xor_i0$15$_i1$15$_o, i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (xor_i0$16$_i1$16$_o, i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (xor_i0$17$_i1$17$_o, i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (xor_i0$18$_i1$18$_o, i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (xor_i0$19$_i1$19$_o, i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (xor_i0$20$_i1$20$_o, i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (xor_i0$21$_i1$21$_o, i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (xor_i0$22$_i1$22$_o, i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (xor_i0$23$_i1$23$_o, i0[23], i1[23]);
  xor \xor_i0[24]_i1[24]  (xor_i0$24$_i1$24$_o, i0[24], i1[24]);
  xor \xor_i0[25]_i1[25]  (xor_i0$25$_i1$25$_o, i0[25], i1[25]);
  xor \xor_i0[26]_i1[26]  (xor_i0$26$_i1$26$_o, i0[26], i1[26]);
  xor \xor_i0[27]_i1[27]  (xor_i0$27$_i1$27$_o, i0[27], i1[27]);
  xor \xor_i0[28]_i1[28]  (xor_i0$28$_i1$28$_o, i0[28], i1[28]);
  xor \xor_i0[29]_i1[29]  (xor_i0$29$_i1$29$_o, i0[29], i1[29]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (xor_i0$3$_i1$3$_o, i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (xor_i0$4$_i1$4$_o, i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (xor_i0$5$_i1$5$_o, i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (xor_i0$6$_i1$6$_o, i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (xor_i0$7$_i1$7$_o, i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (xor_i0$8$_i1$8$_o, i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (xor_i0$9$_i1$9$_o, i0[9], i1[9]);

endmodule 

module binary_mux_s1_w1
  (
  i0,
  i1,
  sel,
  o
  );

  input i0;
  input i1;
  input sel;
  output o;


  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel),
    .o(o));

endmodule 

module ne_w2
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output o;

  wire [1:0] diff;

  or any_diff (o, diff[0], diff[1]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module add_pu30_pu30_o30
  (
  i0,
  i1,
  o
  );

  input [29:0] i0;
  input [29:0] i1;
  output [29:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module add_pu32_pu32_o32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output [31:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module add_pu64_pu64_o64
  (
  i0,
  i1,
  o
  );

  input [63:0] i0;
  input [63:0] i1;
  output [63:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a32;
  wire net_a33;
  wire net_a34;
  wire net_a35;
  wire net_a36;
  wire net_a37;
  wire net_a38;
  wire net_a39;
  wire net_a4;
  wire net_a40;
  wire net_a41;
  wire net_a42;
  wire net_a43;
  wire net_a44;
  wire net_a45;
  wire net_a46;
  wire net_a47;
  wire net_a48;
  wire net_a49;
  wire net_a5;
  wire net_a50;
  wire net_a51;
  wire net_a52;
  wire net_a53;
  wire net_a54;
  wire net_a55;
  wire net_a56;
  wire net_a57;
  wire net_a58;
  wire net_a59;
  wire net_a6;
  wire net_a60;
  wire net_a61;
  wire net_a62;
  wire net_a63;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b32;
  wire net_b33;
  wire net_b34;
  wire net_b35;
  wire net_b36;
  wire net_b37;
  wire net_b38;
  wire net_b39;
  wire net_b4;
  wire net_b40;
  wire net_b41;
  wire net_b42;
  wire net_b43;
  wire net_b44;
  wire net_b45;
  wire net_b46;
  wire net_b47;
  wire net_b48;
  wire net_b49;
  wire net_b5;
  wire net_b50;
  wire net_b51;
  wire net_b52;
  wire net_b53;
  wire net_b54;
  wire net_b55;
  wire net_b56;
  wire net_b57;
  wire net_b58;
  wire net_b59;
  wire net_b6;
  wire net_b60;
  wire net_b61;
  wire net_b62;
  wire net_b63;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout32;
  wire net_cout33;
  wire net_cout34;
  wire net_cout35;
  wire net_cout36;
  wire net_cout37;
  wire net_cout38;
  wire net_cout39;
  wire net_cout4;
  wire net_cout40;
  wire net_cout41;
  wire net_cout42;
  wire net_cout43;
  wire net_cout44;
  wire net_cout45;
  wire net_cout46;
  wire net_cout47;
  wire net_cout48;
  wire net_cout49;
  wire net_cout5;
  wire net_cout50;
  wire net_cout51;
  wire net_cout52;
  wire net_cout53;
  wire net_cout54;
  wire net_cout55;
  wire net_cout56;
  wire net_cout57;
  wire net_cout58;
  wire net_cout59;
  wire net_cout6;
  wire net_cout60;
  wire net_cout61;
  wire net_cout62;
  wire net_cout63;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum32;
  wire net_sum33;
  wire net_sum34;
  wire net_sum35;
  wire net_sum36;
  wire net_sum37;
  wire net_sum38;
  wire net_sum39;
  wire net_sum4;
  wire net_sum40;
  wire net_sum41;
  wire net_sum42;
  wire net_sum43;
  wire net_sum44;
  wire net_sum45;
  wire net_sum46;
  wire net_sum47;
  wire net_sum48;
  wire net_sum49;
  wire net_sum5;
  wire net_sum50;
  wire net_sum51;
  wire net_sum52;
  wire net_sum53;
  wire net_sum54;
  wire net_sum55;
  wire net_sum56;
  wire net_sum57;
  wire net_sum58;
  wire net_sum59;
  wire net_sum6;
  wire net_sum60;
  wire net_sum61;
  wire net_sum62;
  wire net_sum63;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a63 = i0[63];
  assign net_a62 = i0[62];
  assign net_a61 = i0[61];
  assign net_a60 = i0[60];
  assign net_a59 = i0[59];
  assign net_a58 = i0[58];
  assign net_a57 = i0[57];
  assign net_a56 = i0[56];
  assign net_a55 = i0[55];
  assign net_a54 = i0[54];
  assign net_a53 = i0[53];
  assign net_a52 = i0[52];
  assign net_a51 = i0[51];
  assign net_a50 = i0[50];
  assign net_a49 = i0[49];
  assign net_a48 = i0[48];
  assign net_a47 = i0[47];
  assign net_a46 = i0[46];
  assign net_a45 = i0[45];
  assign net_a44 = i0[44];
  assign net_a43 = i0[43];
  assign net_a42 = i0[42];
  assign net_a41 = i0[41];
  assign net_a40 = i0[40];
  assign net_a39 = i0[39];
  assign net_a38 = i0[38];
  assign net_a37 = i0[37];
  assign net_a36 = i0[36];
  assign net_a35 = i0[35];
  assign net_a34 = i0[34];
  assign net_a33 = i0[33];
  assign net_a32 = i0[32];
  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b63 = i1[63];
  assign net_b62 = i1[62];
  assign net_b61 = i1[61];
  assign net_b60 = i1[60];
  assign net_b59 = i1[59];
  assign net_b58 = i1[58];
  assign net_b57 = i1[57];
  assign net_b56 = i1[56];
  assign net_b55 = i1[55];
  assign net_b54 = i1[54];
  assign net_b53 = i1[53];
  assign net_b52 = i1[52];
  assign net_b51 = i1[51];
  assign net_b50 = i1[50];
  assign net_b49 = i1[49];
  assign net_b48 = i1[48];
  assign net_b47 = i1[47];
  assign net_b46 = i1[46];
  assign net_b45 = i1[45];
  assign net_b44 = i1[44];
  assign net_b43 = i1[43];
  assign net_b42 = i1[42];
  assign net_b41 = i1[41];
  assign net_b40 = i1[40];
  assign net_b39 = i1[39];
  assign net_b38 = i1[38];
  assign net_b37 = i1[37];
  assign net_b36 = i1[36];
  assign net_b35 = i1[35];
  assign net_b34 = i1[34];
  assign net_b33 = i1[33];
  assign net_b32 = i1[32];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[63] = net_sum63;
  assign o[62] = net_sum62;
  assign o[61] = net_sum61;
  assign o[60] = net_sum60;
  assign o[59] = net_sum59;
  assign o[58] = net_sum58;
  assign o[57] = net_sum57;
  assign o[56] = net_sum56;
  assign o[55] = net_sum55;
  assign o[54] = net_sum54;
  assign o[53] = net_sum53;
  assign o[52] = net_sum52;
  assign o[51] = net_sum51;
  assign o[50] = net_sum50;
  assign o[49] = net_sum49;
  assign o[48] = net_sum48;
  assign o[47] = net_sum47;
  assign o[46] = net_sum46;
  assign o[45] = net_sum45;
  assign o[44] = net_sum44;
  assign o[43] = net_sum43;
  assign o[42] = net_sum42;
  assign o[41] = net_sum41;
  assign o[40] = net_sum40;
  assign o[39] = net_sum39;
  assign o[38] = net_sum38;
  assign o[37] = net_sum37;
  assign o[36] = net_sum36;
  assign o[35] = net_sum35;
  assign o[34] = net_sum34;
  assign o[33] = net_sum33;
  assign o[32] = net_sum32;
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_32 (
    .a(net_a32),
    .b(net_b32),
    .c(net_cout31),
    .cout(net_cout32),
    .sum(net_sum32));
  AL_FADD comp_33 (
    .a(net_a33),
    .b(net_b33),
    .c(net_cout32),
    .cout(net_cout33),
    .sum(net_sum33));
  AL_FADD comp_34 (
    .a(net_a34),
    .b(net_b34),
    .c(net_cout33),
    .cout(net_cout34),
    .sum(net_sum34));
  AL_FADD comp_35 (
    .a(net_a35),
    .b(net_b35),
    .c(net_cout34),
    .cout(net_cout35),
    .sum(net_sum35));
  AL_FADD comp_36 (
    .a(net_a36),
    .b(net_b36),
    .c(net_cout35),
    .cout(net_cout36),
    .sum(net_sum36));
  AL_FADD comp_37 (
    .a(net_a37),
    .b(net_b37),
    .c(net_cout36),
    .cout(net_cout37),
    .sum(net_sum37));
  AL_FADD comp_38 (
    .a(net_a38),
    .b(net_b38),
    .c(net_cout37),
    .cout(net_cout38),
    .sum(net_sum38));
  AL_FADD comp_39 (
    .a(net_a39),
    .b(net_b39),
    .c(net_cout38),
    .cout(net_cout39),
    .sum(net_sum39));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_40 (
    .a(net_a40),
    .b(net_b40),
    .c(net_cout39),
    .cout(net_cout40),
    .sum(net_sum40));
  AL_FADD comp_41 (
    .a(net_a41),
    .b(net_b41),
    .c(net_cout40),
    .cout(net_cout41),
    .sum(net_sum41));
  AL_FADD comp_42 (
    .a(net_a42),
    .b(net_b42),
    .c(net_cout41),
    .cout(net_cout42),
    .sum(net_sum42));
  AL_FADD comp_43 (
    .a(net_a43),
    .b(net_b43),
    .c(net_cout42),
    .cout(net_cout43),
    .sum(net_sum43));
  AL_FADD comp_44 (
    .a(net_a44),
    .b(net_b44),
    .c(net_cout43),
    .cout(net_cout44),
    .sum(net_sum44));
  AL_FADD comp_45 (
    .a(net_a45),
    .b(net_b45),
    .c(net_cout44),
    .cout(net_cout45),
    .sum(net_sum45));
  AL_FADD comp_46 (
    .a(net_a46),
    .b(net_b46),
    .c(net_cout45),
    .cout(net_cout46),
    .sum(net_sum46));
  AL_FADD comp_47 (
    .a(net_a47),
    .b(net_b47),
    .c(net_cout46),
    .cout(net_cout47),
    .sum(net_sum47));
  AL_FADD comp_48 (
    .a(net_a48),
    .b(net_b48),
    .c(net_cout47),
    .cout(net_cout48),
    .sum(net_sum48));
  AL_FADD comp_49 (
    .a(net_a49),
    .b(net_b49),
    .c(net_cout48),
    .cout(net_cout49),
    .sum(net_sum49));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_50 (
    .a(net_a50),
    .b(net_b50),
    .c(net_cout49),
    .cout(net_cout50),
    .sum(net_sum50));
  AL_FADD comp_51 (
    .a(net_a51),
    .b(net_b51),
    .c(net_cout50),
    .cout(net_cout51),
    .sum(net_sum51));
  AL_FADD comp_52 (
    .a(net_a52),
    .b(net_b52),
    .c(net_cout51),
    .cout(net_cout52),
    .sum(net_sum52));
  AL_FADD comp_53 (
    .a(net_a53),
    .b(net_b53),
    .c(net_cout52),
    .cout(net_cout53),
    .sum(net_sum53));
  AL_FADD comp_54 (
    .a(net_a54),
    .b(net_b54),
    .c(net_cout53),
    .cout(net_cout54),
    .sum(net_sum54));
  AL_FADD comp_55 (
    .a(net_a55),
    .b(net_b55),
    .c(net_cout54),
    .cout(net_cout55),
    .sum(net_sum55));
  AL_FADD comp_56 (
    .a(net_a56),
    .b(net_b56),
    .c(net_cout55),
    .cout(net_cout56),
    .sum(net_sum56));
  AL_FADD comp_57 (
    .a(net_a57),
    .b(net_b57),
    .c(net_cout56),
    .cout(net_cout57),
    .sum(net_sum57));
  AL_FADD comp_58 (
    .a(net_a58),
    .b(net_b58),
    .c(net_cout57),
    .cout(net_cout58),
    .sum(net_sum58));
  AL_FADD comp_59 (
    .a(net_a59),
    .b(net_b59),
    .c(net_cout58),
    .cout(net_cout59),
    .sum(net_sum59));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_60 (
    .a(net_a60),
    .b(net_b60),
    .c(net_cout59),
    .cout(net_cout60),
    .sum(net_sum60));
  AL_FADD comp_61 (
    .a(net_a61),
    .b(net_b61),
    .c(net_cout60),
    .cout(net_cout61),
    .sum(net_sum61));
  AL_FADD comp_62 (
    .a(net_a62),
    .b(net_b62),
    .c(net_cout61),
    .cout(net_cout62),
    .sum(net_sum62));
  AL_FADD comp_63 (
    .a(net_a63),
    .b(net_b63),
    .c(net_cout62),
    .cout(net_cout63),
    .sum(net_sum63));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module reg_ar_ss_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire setout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(setout),
    .reset(reset),
    .set(1'b0),
    .q(q));
  AL_MUX u_set0 (
    .i0(enout),
    .i1(1'b1),
    .sel(set),
    .o(setout));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module eq_w3
  (
  i0,
  i1,
  o
  );

  input [2:0] i0;
  input [2:0] i1;
  output o;

  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$1$_i1$1$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$2$_i1$2$_o;

  not none_diff (o, or_xor_i0$0$_i1$0$_o_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, or_xor_i0$1$_i1$1$_o_o);
  or or_xor_i0$1$_i1$1$_o (or_xor_i0$1$_i1$1$_o_o, xor_i0$1$_i1$1$_o, xor_i0$2$_i1$2$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);

endmodule 

module eq_w1
  (
  i0,
  i1,
  o
  );

  input i0;
  input i1;
  output o;

  wire xor_i0_i1_o;

  not none_diff (o, xor_i0_i1_o);
  xor xor_i0_i1 (xor_i0_i1_o, i0, i1);

endmodule 

module eq_w5
  (
  i0,
  i1,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  output o;

  wire or_or_xor_i0$0$_i1$0_o;
  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$2$_i1$2$_o_o;
  wire or_xor_i0$3$_i1$3$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$2$_i1$2$_o;
  wire xor_i0$3$_i1$3$_o;
  wire xor_i0$4$_i1$4$_o;

  not none_diff (o, or_or_xor_i0$0$_i1$0_o);
  or or_or_xor_i0$0$_i1$0 (or_or_xor_i0$0$_i1$0_o, or_xor_i0$0$_i1$0$_o_o, or_xor_i0$2$_i1$2$_o_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, xor_i0$1$_i1$1$_o);
  or or_xor_i0$2$_i1$2$_o (or_xor_i0$2$_i1$2$_o_o, xor_i0$2$_i1$2$_o, or_xor_i0$3$_i1$3$_o_o);
  or or_xor_i0$3$_i1$3$_o (or_xor_i0$3$_i1$3$_o_o, xor_i0$3$_i1$3$_o, xor_i0$4$_i1$4$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (xor_i0$3$_i1$3$_o, i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (xor_i0$4$_i1$4$_o, i0[4], i1[4]);

endmodule 

module eq_w7
  (
  i0,
  i1,
  o
  );

  input [6:0] i0;
  input [6:0] i1;
  output o;

  wire or_or_xor_i0$0$_i1$0_o;
  wire or_or_xor_i0$3$_i1$3_o;
  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$1$_i1$1$_o_o;
  wire or_xor_i0$3$_i1$3$_o_o;
  wire or_xor_i0$5$_i1$5$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$2$_i1$2$_o;
  wire xor_i0$3$_i1$3$_o;
  wire xor_i0$4$_i1$4$_o;
  wire xor_i0$5$_i1$5$_o;
  wire xor_i0$6$_i1$6$_o;

  not none_diff (o, or_or_xor_i0$0$_i1$0_o);
  or or_or_xor_i0$0$_i1$0 (or_or_xor_i0$0$_i1$0_o, or_xor_i0$0$_i1$0$_o_o, or_or_xor_i0$3$_i1$3_o);
  or or_or_xor_i0$3$_i1$3 (or_or_xor_i0$3$_i1$3_o, or_xor_i0$3$_i1$3$_o_o, or_xor_i0$5$_i1$5$_o_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, or_xor_i0$1$_i1$1$_o_o);
  or or_xor_i0$1$_i1$1$_o (or_xor_i0$1$_i1$1$_o_o, xor_i0$1$_i1$1$_o, xor_i0$2$_i1$2$_o);
  or or_xor_i0$3$_i1$3$_o (or_xor_i0$3$_i1$3$_o_o, xor_i0$3$_i1$3$_o, xor_i0$4$_i1$4$_o);
  or or_xor_i0$5$_i1$5$_o (or_xor_i0$5$_i1$5$_o_o, xor_i0$5$_i1$5$_o, xor_i0$6$_i1$6$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (xor_i0$3$_i1$3$_o, i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (xor_i0$4$_i1$4$_o, i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (xor_i0$5$_i1$5$_o, i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (xor_i0$6$_i1$6$_o, i0[6], i1[6]);

endmodule 

module eq_w32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output o;

  wire or_or_or_or_or_xor_i_o;
  wire or_or_or_or_xor_i0$0_o;
  wire or_or_or_or_xor_i0$1_o;
  wire or_or_or_xor_i0$0$_i_o;
  wire or_or_or_xor_i0$16$__o;
  wire or_or_or_xor_i0$24$__o;
  wire or_or_or_xor_i0$8$_i_o;
  wire or_or_xor_i0$0$_i1$0_o;
  wire or_or_xor_i0$12$_i1$_o;
  wire or_or_xor_i0$16$_i1$_o;
  wire or_or_xor_i0$20$_i1$_o;
  wire or_or_xor_i0$24$_i1$_o;
  wire or_or_xor_i0$28$_i1$_o;
  wire or_or_xor_i0$4$_i1$4_o;
  wire or_or_xor_i0$8$_i1$8_o;
  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$10$_i1$10$_o;
  wire or_xor_i0$12$_i1$12$_o;
  wire or_xor_i0$14$_i1$14$_o;
  wire or_xor_i0$16$_i1$16$_o;
  wire or_xor_i0$18$_i1$18$_o;
  wire or_xor_i0$2$_i1$2$_o_o;
  wire or_xor_i0$20$_i1$20$_o;
  wire or_xor_i0$22$_i1$22$_o;
  wire or_xor_i0$24$_i1$24$_o;
  wire or_xor_i0$26$_i1$26$_o;
  wire or_xor_i0$28$_i1$28$_o;
  wire or_xor_i0$30$_i1$30$_o;
  wire or_xor_i0$4$_i1$4$_o_o;
  wire or_xor_i0$6$_i1$6$_o_o;
  wire or_xor_i0$8$_i1$8$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$10$_i1$10$_o;
  wire xor_i0$11$_i1$11$_o;
  wire xor_i0$12$_i1$12$_o;
  wire xor_i0$13$_i1$13$_o;
  wire xor_i0$14$_i1$14$_o;
  wire xor_i0$15$_i1$15$_o;
  wire xor_i0$16$_i1$16$_o;
  wire xor_i0$17$_i1$17$_o;
  wire xor_i0$18$_i1$18$_o;
  wire xor_i0$19$_i1$19$_o;
  wire xor_i0$2$_i1$2$_o;
  wire xor_i0$20$_i1$20$_o;
  wire xor_i0$21$_i1$21$_o;
  wire xor_i0$22$_i1$22$_o;
  wire xor_i0$23$_i1$23$_o;
  wire xor_i0$24$_i1$24$_o;
  wire xor_i0$25$_i1$25$_o;
  wire xor_i0$26$_i1$26$_o;
  wire xor_i0$27$_i1$27$_o;
  wire xor_i0$28$_i1$28$_o;
  wire xor_i0$29$_i1$29$_o;
  wire xor_i0$3$_i1$3$_o;
  wire xor_i0$30$_i1$30$_o;
  wire xor_i0$31$_i1$31$_o;
  wire xor_i0$4$_i1$4$_o;
  wire xor_i0$5$_i1$5$_o;
  wire xor_i0$6$_i1$6$_o;
  wire xor_i0$7$_i1$7$_o;
  wire xor_i0$8$_i1$8$_o;
  wire xor_i0$9$_i1$9$_o;

  not none_diff (o, or_or_or_or_or_xor_i_o);
  or or_or_or_or_or_xor_i (or_or_or_or_or_xor_i_o, or_or_or_or_xor_i0$0_o, or_or_or_or_xor_i0$1_o);
  or or_or_or_or_xor_i0$0 (or_or_or_or_xor_i0$0_o, or_or_or_xor_i0$0$_i_o, or_or_or_xor_i0$8$_i_o);
  or or_or_or_or_xor_i0$1 (or_or_or_or_xor_i0$1_o, or_or_or_xor_i0$16$__o, or_or_or_xor_i0$24$__o);
  or or_or_or_xor_i0$0$_i (or_or_or_xor_i0$0$_i_o, or_or_xor_i0$0$_i1$0_o, or_or_xor_i0$4$_i1$4_o);
  or or_or_or_xor_i0$16$_ (or_or_or_xor_i0$16$__o, or_or_xor_i0$16$_i1$_o, or_or_xor_i0$20$_i1$_o);
  or or_or_or_xor_i0$24$_ (or_or_or_xor_i0$24$__o, or_or_xor_i0$24$_i1$_o, or_or_xor_i0$28$_i1$_o);
  or or_or_or_xor_i0$8$_i (or_or_or_xor_i0$8$_i_o, or_or_xor_i0$8$_i1$8_o, or_or_xor_i0$12$_i1$_o);
  or or_or_xor_i0$0$_i1$0 (or_or_xor_i0$0$_i1$0_o, or_xor_i0$0$_i1$0$_o_o, or_xor_i0$2$_i1$2$_o_o);
  or or_or_xor_i0$12$_i1$ (or_or_xor_i0$12$_i1$_o, or_xor_i0$12$_i1$12$_o, or_xor_i0$14$_i1$14$_o);
  or or_or_xor_i0$16$_i1$ (or_or_xor_i0$16$_i1$_o, or_xor_i0$16$_i1$16$_o, or_xor_i0$18$_i1$18$_o);
  or or_or_xor_i0$20$_i1$ (or_or_xor_i0$20$_i1$_o, or_xor_i0$20$_i1$20$_o, or_xor_i0$22$_i1$22$_o);
  or or_or_xor_i0$24$_i1$ (or_or_xor_i0$24$_i1$_o, or_xor_i0$24$_i1$24$_o, or_xor_i0$26$_i1$26$_o);
  or or_or_xor_i0$28$_i1$ (or_or_xor_i0$28$_i1$_o, or_xor_i0$28$_i1$28$_o, or_xor_i0$30$_i1$30$_o);
  or or_or_xor_i0$4$_i1$4 (or_or_xor_i0$4$_i1$4_o, or_xor_i0$4$_i1$4$_o_o, or_xor_i0$6$_i1$6$_o_o);
  or or_or_xor_i0$8$_i1$8 (or_or_xor_i0$8$_i1$8_o, or_xor_i0$8$_i1$8$_o_o, or_xor_i0$10$_i1$10$_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, xor_i0$1$_i1$1$_o);
  or or_xor_i0$10$_i1$10$ (or_xor_i0$10$_i1$10$_o, xor_i0$10$_i1$10$_o, xor_i0$11$_i1$11$_o);
  or or_xor_i0$12$_i1$12$ (or_xor_i0$12$_i1$12$_o, xor_i0$12$_i1$12$_o, xor_i0$13$_i1$13$_o);
  or or_xor_i0$14$_i1$14$ (or_xor_i0$14$_i1$14$_o, xor_i0$14$_i1$14$_o, xor_i0$15$_i1$15$_o);
  or or_xor_i0$16$_i1$16$ (or_xor_i0$16$_i1$16$_o, xor_i0$16$_i1$16$_o, xor_i0$17$_i1$17$_o);
  or or_xor_i0$18$_i1$18$ (or_xor_i0$18$_i1$18$_o, xor_i0$18$_i1$18$_o, xor_i0$19$_i1$19$_o);
  or or_xor_i0$2$_i1$2$_o (or_xor_i0$2$_i1$2$_o_o, xor_i0$2$_i1$2$_o, xor_i0$3$_i1$3$_o);
  or or_xor_i0$20$_i1$20$ (or_xor_i0$20$_i1$20$_o, xor_i0$20$_i1$20$_o, xor_i0$21$_i1$21$_o);
  or or_xor_i0$22$_i1$22$ (or_xor_i0$22$_i1$22$_o, xor_i0$22$_i1$22$_o, xor_i0$23$_i1$23$_o);
  or or_xor_i0$24$_i1$24$ (or_xor_i0$24$_i1$24$_o, xor_i0$24$_i1$24$_o, xor_i0$25$_i1$25$_o);
  or or_xor_i0$26$_i1$26$ (or_xor_i0$26$_i1$26$_o, xor_i0$26$_i1$26$_o, xor_i0$27$_i1$27$_o);
  or or_xor_i0$28$_i1$28$ (or_xor_i0$28$_i1$28$_o, xor_i0$28$_i1$28$_o, xor_i0$29$_i1$29$_o);
  or or_xor_i0$30$_i1$30$ (or_xor_i0$30$_i1$30$_o, xor_i0$30$_i1$30$_o, xor_i0$31$_i1$31$_o);
  or or_xor_i0$4$_i1$4$_o (or_xor_i0$4$_i1$4$_o_o, xor_i0$4$_i1$4$_o, xor_i0$5$_i1$5$_o);
  or or_xor_i0$6$_i1$6$_o (or_xor_i0$6$_i1$6$_o_o, xor_i0$6$_i1$6$_o, xor_i0$7$_i1$7$_o);
  or or_xor_i0$8$_i1$8$_o (or_xor_i0$8$_i1$8$_o_o, xor_i0$8$_i1$8$_o, xor_i0$9$_i1$9$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (xor_i0$10$_i1$10$_o, i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (xor_i0$11$_i1$11$_o, i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (xor_i0$12$_i1$12$_o, i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (xor_i0$13$_i1$13$_o, i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (xor_i0$14$_i1$14$_o, i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (xor_i0$15$_i1$15$_o, i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (xor_i0$16$_i1$16$_o, i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (xor_i0$17$_i1$17$_o, i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (xor_i0$18$_i1$18$_o, i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (xor_i0$19$_i1$19$_o, i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (xor_i0$20$_i1$20$_o, i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (xor_i0$21$_i1$21$_o, i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (xor_i0$22$_i1$22$_o, i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (xor_i0$23$_i1$23$_o, i0[23], i1[23]);
  xor \xor_i0[24]_i1[24]  (xor_i0$24$_i1$24$_o, i0[24], i1[24]);
  xor \xor_i0[25]_i1[25]  (xor_i0$25$_i1$25$_o, i0[25], i1[25]);
  xor \xor_i0[26]_i1[26]  (xor_i0$26$_i1$26$_o, i0[26], i1[26]);
  xor \xor_i0[27]_i1[27]  (xor_i0$27$_i1$27$_o, i0[27], i1[27]);
  xor \xor_i0[28]_i1[28]  (xor_i0$28$_i1$28$_o, i0[28], i1[28]);
  xor \xor_i0[29]_i1[29]  (xor_i0$29$_i1$29$_o, i0[29], i1[29]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);
  xor \xor_i0[30]_i1[30]  (xor_i0$30$_i1$30$_o, i0[30], i1[30]);
  xor \xor_i0[31]_i1[31]  (xor_i0$31$_i1$31$_o, i0[31], i1[31]);
  xor \xor_i0[3]_i1[3]  (xor_i0$3$_i1$3$_o, i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (xor_i0$4$_i1$4$_o, i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (xor_i0$5$_i1$5$_o, i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (xor_i0$6$_i1$6$_o, i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (xor_i0$7$_i1$7$_o, i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (xor_i0$8$_i1$8$_o, i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (xor_i0$9$_i1$9$_o, i0[9], i1[9]);

endmodule 

module eq_w8
  (
  i0,
  i1,
  o
  );

  input [7:0] i0;
  input [7:0] i1;
  output o;

  wire or_or_or_xor_i0$0$_i_o;
  wire or_or_xor_i0$0$_i1$0_o;
  wire or_or_xor_i0$4$_i1$4_o;
  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$2$_i1$2$_o_o;
  wire or_xor_i0$4$_i1$4$_o_o;
  wire or_xor_i0$6$_i1$6$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$2$_i1$2$_o;
  wire xor_i0$3$_i1$3$_o;
  wire xor_i0$4$_i1$4$_o;
  wire xor_i0$5$_i1$5$_o;
  wire xor_i0$6$_i1$6$_o;
  wire xor_i0$7$_i1$7$_o;

  not none_diff (o, or_or_or_xor_i0$0$_i_o);
  or or_or_or_xor_i0$0$_i (or_or_or_xor_i0$0$_i_o, or_or_xor_i0$0$_i1$0_o, or_or_xor_i0$4$_i1$4_o);
  or or_or_xor_i0$0$_i1$0 (or_or_xor_i0$0$_i1$0_o, or_xor_i0$0$_i1$0$_o_o, or_xor_i0$2$_i1$2$_o_o);
  or or_or_xor_i0$4$_i1$4 (or_or_xor_i0$4$_i1$4_o, or_xor_i0$4$_i1$4$_o_o, or_xor_i0$6$_i1$6$_o_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, xor_i0$1$_i1$1$_o);
  or or_xor_i0$2$_i1$2$_o (or_xor_i0$2$_i1$2$_o_o, xor_i0$2$_i1$2$_o, xor_i0$3$_i1$3$_o);
  or or_xor_i0$4$_i1$4$_o (or_xor_i0$4$_i1$4$_o_o, xor_i0$4$_i1$4$_o, xor_i0$5$_i1$5$_o);
  or or_xor_i0$6$_i1$6$_o (or_xor_i0$6$_i1$6$_o_o, xor_i0$6$_i1$6$_o, xor_i0$7$_i1$7$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (xor_i0$3$_i1$3$_o, i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (xor_i0$4$_i1$4$_o, i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (xor_i0$5$_i1$5$_o, i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (xor_i0$6$_i1$6$_o, i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (xor_i0$7$_i1$7$_o, i0[7], i1[7]);

endmodule 

module lt_u32_u32
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [31:0] i0;
  input [31:0] i1;
  output o;

  wire [31:0] diff;
  wire diff_12_18;
  wire diff_19_26;
  wire diff_27_31;
  wire diff_6_11;
  wire less_12_18;
  wire \less_12_18_inst/diff_0 ;
  wire \less_12_18_inst/diff_1 ;
  wire \less_12_18_inst/diff_2 ;
  wire \less_12_18_inst/diff_3 ;
  wire \less_12_18_inst/diff_4 ;
  wire \less_12_18_inst/diff_5 ;
  wire \less_12_18_inst/diff_6 ;
  wire \less_12_18_inst/o_0 ;
  wire \less_12_18_inst/o_1 ;
  wire \less_12_18_inst/o_2 ;
  wire \less_12_18_inst/o_3 ;
  wire \less_12_18_inst/o_4 ;
  wire \less_12_18_inst/o_5 ;
  wire less_19_26;
  wire \less_19_26_inst/diff_0 ;
  wire \less_19_26_inst/diff_1 ;
  wire \less_19_26_inst/diff_2 ;
  wire \less_19_26_inst/diff_3 ;
  wire \less_19_26_inst/diff_4 ;
  wire \less_19_26_inst/diff_5 ;
  wire \less_19_26_inst/diff_6 ;
  wire \less_19_26_inst/diff_7 ;
  wire \less_19_26_inst/o_0 ;
  wire \less_19_26_inst/o_1 ;
  wire \less_19_26_inst/o_2 ;
  wire \less_19_26_inst/o_3 ;
  wire \less_19_26_inst/o_4 ;
  wire \less_19_26_inst/o_5 ;
  wire \less_19_26_inst/o_6 ;
  wire less_27_31;
  wire \less_27_31_inst/diff_0 ;
  wire \less_27_31_inst/diff_1 ;
  wire \less_27_31_inst/diff_2 ;
  wire \less_27_31_inst/diff_3 ;
  wire \less_27_31_inst/diff_4 ;
  wire \less_27_31_inst/o_0 ;
  wire \less_27_31_inst/o_1 ;
  wire \less_27_31_inst/o_2 ;
  wire \less_27_31_inst/o_3 ;
  wire less_6_11;
  wire \less_6_11_inst/diff_0 ;
  wire \less_6_11_inst/diff_1 ;
  wire \less_6_11_inst/diff_2 ;
  wire \less_6_11_inst/diff_3 ;
  wire \less_6_11_inst/diff_4 ;
  wire \less_6_11_inst/diff_5 ;
  wire \less_6_11_inst/o_0 ;
  wire \less_6_11_inst/o_1 ;
  wire \less_6_11_inst/o_2 ;
  wire \less_6_11_inst/o_3 ;
  wire \less_6_11_inst/o_4 ;
  wire o_0;
  wire o_1;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;
  wire o_6;
  wire o_7;
  wire o_8;

  or any_diff_12_18 (diff_12_18, diff[12], diff[13], diff[14], diff[15], diff[16], diff[17], diff[18]);
  or any_diff_19_26 (diff_19_26, diff[19], diff[20], diff[21], diff[22], diff[23], diff[24], diff[25], diff[26]);
  or any_diff_27_31 (diff_27_31, diff[27], diff[28], diff[29], diff[30], diff[31]);
  or any_diff_6_11 (diff_6_11, diff[6], diff[7], diff[8], diff[9], diff[10], diff[11]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_12 (diff[12], i0[12], i1[12]);
  xor diff_13 (diff[13], i0[13], i1[13]);
  xor diff_14 (diff[14], i0[14], i1[14]);
  xor diff_15 (diff[15], i0[15], i1[15]);
  xor diff_16 (diff[16], i0[16], i1[16]);
  xor diff_17 (diff[17], i0[17], i1[17]);
  xor diff_18 (diff[18], i0[18], i1[18]);
  xor diff_19 (diff[19], i0[19], i1[19]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_20 (diff[20], i0[20], i1[20]);
  xor diff_21 (diff[21], i0[21], i1[21]);
  xor diff_22 (diff[22], i0[22], i1[22]);
  xor diff_23 (diff[23], i0[23], i1[23]);
  xor diff_24 (diff[24], i0[24], i1[24]);
  xor diff_25 (diff[25], i0[25], i1[25]);
  xor diff_26 (diff[26], i0[26], i1[26]);
  xor diff_27 (diff[27], i0[27], i1[27]);
  xor diff_28 (diff[28], i0[28], i1[28]);
  xor diff_29 (diff[29], i0[29], i1[29]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_30 (diff[30], i0[30], i1[30]);
  xor diff_31 (diff[31], i0[31], i1[31]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);
  AL_MUX \less_12_18_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[12]),
    .sel(\less_12_18_inst/diff_0 ),
    .o(\less_12_18_inst/o_0 ));
  AL_MUX \less_12_18_inst/mux_1  (
    .i0(\less_12_18_inst/o_0 ),
    .i1(i1[13]),
    .sel(\less_12_18_inst/diff_1 ),
    .o(\less_12_18_inst/o_1 ));
  AL_MUX \less_12_18_inst/mux_2  (
    .i0(\less_12_18_inst/o_1 ),
    .i1(i1[14]),
    .sel(\less_12_18_inst/diff_2 ),
    .o(\less_12_18_inst/o_2 ));
  AL_MUX \less_12_18_inst/mux_3  (
    .i0(\less_12_18_inst/o_2 ),
    .i1(i1[15]),
    .sel(\less_12_18_inst/diff_3 ),
    .o(\less_12_18_inst/o_3 ));
  AL_MUX \less_12_18_inst/mux_4  (
    .i0(\less_12_18_inst/o_3 ),
    .i1(i1[16]),
    .sel(\less_12_18_inst/diff_4 ),
    .o(\less_12_18_inst/o_4 ));
  AL_MUX \less_12_18_inst/mux_5  (
    .i0(\less_12_18_inst/o_4 ),
    .i1(i1[17]),
    .sel(\less_12_18_inst/diff_5 ),
    .o(\less_12_18_inst/o_5 ));
  AL_MUX \less_12_18_inst/mux_6  (
    .i0(\less_12_18_inst/o_5 ),
    .i1(i1[18]),
    .sel(\less_12_18_inst/diff_6 ),
    .o(less_12_18));
  xor \less_12_18_inst/xor_0  (\less_12_18_inst/diff_0 , i0[12], i1[12]);
  xor \less_12_18_inst/xor_1  (\less_12_18_inst/diff_1 , i0[13], i1[13]);
  xor \less_12_18_inst/xor_2  (\less_12_18_inst/diff_2 , i0[14], i1[14]);
  xor \less_12_18_inst/xor_3  (\less_12_18_inst/diff_3 , i0[15], i1[15]);
  xor \less_12_18_inst/xor_4  (\less_12_18_inst/diff_4 , i0[16], i1[16]);
  xor \less_12_18_inst/xor_5  (\less_12_18_inst/diff_5 , i0[17], i1[17]);
  xor \less_12_18_inst/xor_6  (\less_12_18_inst/diff_6 , i0[18], i1[18]);
  AL_MUX \less_19_26_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[19]),
    .sel(\less_19_26_inst/diff_0 ),
    .o(\less_19_26_inst/o_0 ));
  AL_MUX \less_19_26_inst/mux_1  (
    .i0(\less_19_26_inst/o_0 ),
    .i1(i1[20]),
    .sel(\less_19_26_inst/diff_1 ),
    .o(\less_19_26_inst/o_1 ));
  AL_MUX \less_19_26_inst/mux_2  (
    .i0(\less_19_26_inst/o_1 ),
    .i1(i1[21]),
    .sel(\less_19_26_inst/diff_2 ),
    .o(\less_19_26_inst/o_2 ));
  AL_MUX \less_19_26_inst/mux_3  (
    .i0(\less_19_26_inst/o_2 ),
    .i1(i1[22]),
    .sel(\less_19_26_inst/diff_3 ),
    .o(\less_19_26_inst/o_3 ));
  AL_MUX \less_19_26_inst/mux_4  (
    .i0(\less_19_26_inst/o_3 ),
    .i1(i1[23]),
    .sel(\less_19_26_inst/diff_4 ),
    .o(\less_19_26_inst/o_4 ));
  AL_MUX \less_19_26_inst/mux_5  (
    .i0(\less_19_26_inst/o_4 ),
    .i1(i1[24]),
    .sel(\less_19_26_inst/diff_5 ),
    .o(\less_19_26_inst/o_5 ));
  AL_MUX \less_19_26_inst/mux_6  (
    .i0(\less_19_26_inst/o_5 ),
    .i1(i1[25]),
    .sel(\less_19_26_inst/diff_6 ),
    .o(\less_19_26_inst/o_6 ));
  AL_MUX \less_19_26_inst/mux_7  (
    .i0(\less_19_26_inst/o_6 ),
    .i1(i1[26]),
    .sel(\less_19_26_inst/diff_7 ),
    .o(less_19_26));
  xor \less_19_26_inst/xor_0  (\less_19_26_inst/diff_0 , i0[19], i1[19]);
  xor \less_19_26_inst/xor_1  (\less_19_26_inst/diff_1 , i0[20], i1[20]);
  xor \less_19_26_inst/xor_2  (\less_19_26_inst/diff_2 , i0[21], i1[21]);
  xor \less_19_26_inst/xor_3  (\less_19_26_inst/diff_3 , i0[22], i1[22]);
  xor \less_19_26_inst/xor_4  (\less_19_26_inst/diff_4 , i0[23], i1[23]);
  xor \less_19_26_inst/xor_5  (\less_19_26_inst/diff_5 , i0[24], i1[24]);
  xor \less_19_26_inst/xor_6  (\less_19_26_inst/diff_6 , i0[25], i1[25]);
  xor \less_19_26_inst/xor_7  (\less_19_26_inst/diff_7 , i0[26], i1[26]);
  AL_MUX \less_27_31_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[27]),
    .sel(\less_27_31_inst/diff_0 ),
    .o(\less_27_31_inst/o_0 ));
  AL_MUX \less_27_31_inst/mux_1  (
    .i0(\less_27_31_inst/o_0 ),
    .i1(i1[28]),
    .sel(\less_27_31_inst/diff_1 ),
    .o(\less_27_31_inst/o_1 ));
  AL_MUX \less_27_31_inst/mux_2  (
    .i0(\less_27_31_inst/o_1 ),
    .i1(i1[29]),
    .sel(\less_27_31_inst/diff_2 ),
    .o(\less_27_31_inst/o_2 ));
  AL_MUX \less_27_31_inst/mux_3  (
    .i0(\less_27_31_inst/o_2 ),
    .i1(i1[30]),
    .sel(\less_27_31_inst/diff_3 ),
    .o(\less_27_31_inst/o_3 ));
  AL_MUX \less_27_31_inst/mux_4  (
    .i0(\less_27_31_inst/o_3 ),
    .i1(i1[31]),
    .sel(\less_27_31_inst/diff_4 ),
    .o(less_27_31));
  xor \less_27_31_inst/xor_0  (\less_27_31_inst/diff_0 , i0[27], i1[27]);
  xor \less_27_31_inst/xor_1  (\less_27_31_inst/diff_1 , i0[28], i1[28]);
  xor \less_27_31_inst/xor_2  (\less_27_31_inst/diff_2 , i0[29], i1[29]);
  xor \less_27_31_inst/xor_3  (\less_27_31_inst/diff_3 , i0[30], i1[30]);
  xor \less_27_31_inst/xor_4  (\less_27_31_inst/diff_4 , i0[31], i1[31]);
  AL_MUX \less_6_11_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[6]),
    .sel(\less_6_11_inst/diff_0 ),
    .o(\less_6_11_inst/o_0 ));
  AL_MUX \less_6_11_inst/mux_1  (
    .i0(\less_6_11_inst/o_0 ),
    .i1(i1[7]),
    .sel(\less_6_11_inst/diff_1 ),
    .o(\less_6_11_inst/o_1 ));
  AL_MUX \less_6_11_inst/mux_2  (
    .i0(\less_6_11_inst/o_1 ),
    .i1(i1[8]),
    .sel(\less_6_11_inst/diff_2 ),
    .o(\less_6_11_inst/o_2 ));
  AL_MUX \less_6_11_inst/mux_3  (
    .i0(\less_6_11_inst/o_2 ),
    .i1(i1[9]),
    .sel(\less_6_11_inst/diff_3 ),
    .o(\less_6_11_inst/o_3 ));
  AL_MUX \less_6_11_inst/mux_4  (
    .i0(\less_6_11_inst/o_3 ),
    .i1(i1[10]),
    .sel(\less_6_11_inst/diff_4 ),
    .o(\less_6_11_inst/o_4 ));
  AL_MUX \less_6_11_inst/mux_5  (
    .i0(\less_6_11_inst/o_4 ),
    .i1(i1[11]),
    .sel(\less_6_11_inst/diff_5 ),
    .o(less_6_11));
  xor \less_6_11_inst/xor_0  (\less_6_11_inst/diff_0 , i0[6], i1[6]);
  xor \less_6_11_inst/xor_1  (\less_6_11_inst/diff_1 , i0[7], i1[7]);
  xor \less_6_11_inst/xor_2  (\less_6_11_inst/diff_2 , i0[8], i1[8]);
  xor \less_6_11_inst/xor_3  (\less_6_11_inst/diff_3 , i0[9], i1[9]);
  xor \less_6_11_inst/xor_4  (\less_6_11_inst/diff_4 , i0[10], i1[10]);
  xor \less_6_11_inst/xor_5  (\less_6_11_inst/diff_5 , i0[11], i1[11]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(i1[4]),
    .sel(diff[4]),
    .o(o_4));
  AL_MUX mux_5 (
    .i0(o_4),
    .i1(i1[5]),
    .sel(diff[5]),
    .o(o_5));
  AL_MUX mux_6 (
    .i0(o_5),
    .i1(less_6_11),
    .sel(diff_6_11),
    .o(o_6));
  AL_MUX mux_7 (
    .i0(o_6),
    .i1(less_12_18),
    .sel(diff_12_18),
    .o(o_7));
  AL_MUX mux_8 (
    .i0(o_7),
    .i1(less_19_26),
    .sel(diff_19_26),
    .o(o_8));
  AL_MUX mux_9 (
    .i0(o_8),
    .i1(less_27_31),
    .sel(diff_27_31),
    .o(o));

endmodule 

module lt_u5_u5
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [4:0] i0;
  input [4:0] i1;
  output o;

  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire diff_0;
  wire diff_1;
  wire diff_2;
  wire diff_3;
  wire diff_4;
  wire net_cin;
  wire o_0;
  wire o_1;
  wire o_2;
  wire o_3;
  wire o_4;

  assign net_cin = ci;
  assign a_4 = i0[4];
  assign a_3 = i0[3];
  assign a_2 = i0[2];
  assign a_1 = i0[1];
  assign a_0 = i0[0];
  assign b_4 = i1[4];
  assign b_3 = i1[3];
  assign b_2 = i1[2];
  assign b_1 = i1[1];
  assign b_0 = i1[0];
  assign o = o_4;
  AL_MUX mux_0 (
    .i0(net_cin),
    .i1(b_0),
    .sel(diff_0),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(b_1),
    .sel(diff_1),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(b_2),
    .sel(diff_2),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(b_3),
    .sel(diff_3),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(b_4),
    .sel(diff_4),
    .o(o_4));
  xor xor_0 (diff_0, a_0, b_0);
  xor xor_1 (diff_1, a_1, b_1);
  xor xor_2 (diff_2, a_2, b_2);
  xor xor_3 (diff_3, a_3, b_3);
  xor xor_4 (diff_4, a_4, b_4);

endmodule 

module binary_mux_s2_w1
  (
  i0,
  i1,
  i2,
  i3,
  sel,
  o
  );

  input i0;
  input i1;
  input i2;
  input i3;
  input [1:0] sel;
  output o;

  wire  B0_0;
  wire  B0_1;

  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel[0]),
    .o(B0_0));
  AL_MUX al_mux_b0_0_1 (
    .i0(i2),
    .i1(i3),
    .sel(sel[0]),
    .o(B0_1));
  AL_MUX al_mux_b0_1_0 (
    .i0(B0_0),
    .i1(B0_1),
    .sel(sel[1]),
    .o(o));

endmodule 

module binary_mux_s3_w1
  (
  i0,
  i1,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  sel,
  o
  );

  input i0;
  input i1;
  input i2;
  input i3;
  input i4;
  input i5;
  input i6;
  input i7;
  input [2:0] sel;
  output o;

  wire  B0_0;
  wire  B0_1;
  wire  B0_2;
  wire  B0_3;
  wire  B1_0;
  wire  B1_1;

  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel[0]),
    .o(B0_0));
  AL_MUX al_mux_b0_0_1 (
    .i0(i2),
    .i1(i3),
    .sel(sel[0]),
    .o(B0_1));
  AL_MUX al_mux_b0_0_2 (
    .i0(i4),
    .i1(i5),
    .sel(sel[0]),
    .o(B0_2));
  AL_MUX al_mux_b0_0_3 (
    .i0(i6),
    .i1(i7),
    .sel(sel[0]),
    .o(B0_3));
  AL_MUX al_mux_b0_1_0 (
    .i0(B0_0),
    .i1(B0_1),
    .sel(sel[1]),
    .o(B1_0));
  AL_MUX al_mux_b0_1_1 (
    .i0(B0_2),
    .i1(B0_3),
    .sel(sel[1]),
    .o(B1_1));
  AL_MUX al_mux_b0_2_0 (
    .i0(B1_0),
    .i1(B1_1),
    .sel(sel[2]),
    .o(o));

endmodule 

module ne_w5
  (
  i0,
  i1,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  output o;

  wire [4:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2], diff[3], diff[4]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);

endmodule 

module ne_w1
  (
  i0,
  i1,
  o
  );

  input i0;
  input i1;
  output o;


  xor diff_0 (o, i0, i1);

endmodule 

module reg_sr_ss_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;
  wire setout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(setout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(1'b0),
    .q(q));
  AL_MUX u_set0 (
    .i0(enout),
    .i1(1'b1),
    .sel(set),
    .o(setout));

endmodule 

module add_pu32_mu32_o32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output [31:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb10;
  wire net_nb11;
  wire net_nb12;
  wire net_nb13;
  wire net_nb14;
  wire net_nb15;
  wire net_nb16;
  wire net_nb17;
  wire net_nb18;
  wire net_nb19;
  wire net_nb2;
  wire net_nb20;
  wire net_nb21;
  wire net_nb22;
  wire net_nb23;
  wire net_nb24;
  wire net_nb25;
  wire net_nb26;
  wire net_nb27;
  wire net_nb28;
  wire net_nb29;
  wire net_nb3;
  wire net_nb30;
  wire net_nb31;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_nb10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_nb11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_nb12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_nb13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_nb14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_nb15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_nb16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_nb17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_nb18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_nb19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_nb20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_nb21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_nb22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_nb23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_nb24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_nb25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_nb26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_nb27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_nb28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_nb29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_nb30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_nb31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b10 (net_nb10, net_b10);
  not inv_b11 (net_nb11, net_b11);
  not inv_b12 (net_nb12, net_b12);
  not inv_b13 (net_nb13, net_b13);
  not inv_b14 (net_nb14, net_b14);
  not inv_b15 (net_nb15, net_b15);
  not inv_b16 (net_nb16, net_b16);
  not inv_b17 (net_nb17, net_b17);
  not inv_b18 (net_nb18, net_b18);
  not inv_b19 (net_nb19, net_b19);
  not inv_b2 (net_nb2, net_b2);
  not inv_b20 (net_nb20, net_b20);
  not inv_b21 (net_nb21, net_b21);
  not inv_b22 (net_nb22, net_b22);
  not inv_b23 (net_nb23, net_b23);
  not inv_b24 (net_nb24, net_b24);
  not inv_b25 (net_nb25, net_b25);
  not inv_b26 (net_nb26, net_b26);
  not inv_b27 (net_nb27, net_b27);
  not inv_b28 (net_nb28, net_b28);
  not inv_b29 (net_nb29, net_b29);
  not inv_b3 (net_nb3, net_b3);
  not inv_b30 (net_nb30, net_b30);
  not inv_b31 (net_nb31, net_b31);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);

endmodule 

module add_pu5_mu5_o5
  (
  i0,
  i1,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  output [4:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_nb0;
  wire net_nb1;
  wire net_nb2;
  wire net_nb3;
  wire net_nb4;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;

  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);

endmodule 

module add_pu4_pu4_o4
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output [3:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;

  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));

endmodule 

module eq_w4
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output o;

  wire or_or_xor_i0$0$_i1$0_o;
  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$2$_i1$2$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$2$_i1$2$_o;
  wire xor_i0$3$_i1$3$_o;

  not none_diff (o, or_or_xor_i0$0$_i1$0_o);
  or or_or_xor_i0$0$_i1$0 (or_or_xor_i0$0$_i1$0_o, or_xor_i0$0$_i1$0$_o_o, or_xor_i0$2$_i1$2$_o_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, xor_i0$1$_i1$1$_o);
  or or_xor_i0$2$_i1$2$_o (or_xor_i0$2$_i1$2$_o_o, xor_i0$2$_i1$2$_o, xor_i0$3$_i1$3$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (xor_i0$3$_i1$3$_o, i0[3], i1[3]);

endmodule 

module lt_u4_u4
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [3:0] i0;
  input [3:0] i1;
  output o;

  wire [3:0] diff;
  wire o_0;
  wire o_1;
  wire o_2;

  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o));

endmodule 

module binary_mux_s4_w1
  (
  i0,
  i1,
  i10,
  i11,
  i12,
  i13,
  i14,
  i15,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  sel,
  o
  );

  input i0;
  input i1;
  input i10;
  input i11;
  input i12;
  input i13;
  input i14;
  input i15;
  input i2;
  input i3;
  input i4;
  input i5;
  input i6;
  input i7;
  input i8;
  input i9;
  input [3:0] sel;
  output o;

  wire  B0_0;
  wire  B0_1;
  wire  B0_2;
  wire  B0_3;
  wire  B0_4;
  wire  B0_5;
  wire  B0_6;
  wire  B0_7;
  wire  B1_0;
  wire  B1_1;
  wire  B1_2;
  wire  B1_3;
  wire  B2_0;
  wire  B2_1;

  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel[0]),
    .o(B0_0));
  AL_MUX al_mux_b0_0_1 (
    .i0(i2),
    .i1(i3),
    .sel(sel[0]),
    .o(B0_1));
  AL_MUX al_mux_b0_0_2 (
    .i0(i4),
    .i1(i5),
    .sel(sel[0]),
    .o(B0_2));
  AL_MUX al_mux_b0_0_3 (
    .i0(i6),
    .i1(i7),
    .sel(sel[0]),
    .o(B0_3));
  AL_MUX al_mux_b0_0_4 (
    .i0(i8),
    .i1(i9),
    .sel(sel[0]),
    .o(B0_4));
  AL_MUX al_mux_b0_0_5 (
    .i0(i10),
    .i1(i11),
    .sel(sel[0]),
    .o(B0_5));
  AL_MUX al_mux_b0_0_6 (
    .i0(i12),
    .i1(i13),
    .sel(sel[0]),
    .o(B0_6));
  AL_MUX al_mux_b0_0_7 (
    .i0(i14),
    .i1(i15),
    .sel(sel[0]),
    .o(B0_7));
  AL_MUX al_mux_b0_1_0 (
    .i0(B0_0),
    .i1(B0_1),
    .sel(sel[1]),
    .o(B1_0));
  AL_MUX al_mux_b0_1_1 (
    .i0(B0_2),
    .i1(B0_3),
    .sel(sel[1]),
    .o(B1_1));
  AL_MUX al_mux_b0_1_2 (
    .i0(B0_4),
    .i1(B0_5),
    .sel(sel[1]),
    .o(B1_2));
  AL_MUX al_mux_b0_1_3 (
    .i0(B0_6),
    .i1(B0_7),
    .sel(sel[1]),
    .o(B1_3));
  AL_MUX al_mux_b0_2_0 (
    .i0(B1_0),
    .i1(B1_1),
    .sel(sel[2]),
    .o(B2_0));
  AL_MUX al_mux_b0_2_1 (
    .i0(B1_2),
    .i1(B1_3),
    .sel(sel[2]),
    .o(B2_1));
  AL_MUX al_mux_b0_3_0 (
    .i0(B2_0),
    .i1(B2_1),
    .sel(sel[3]),
    .o(o));

endmodule 

module ne_w4
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output o;

  wire [3:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2], diff[3]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);

endmodule 

module add_pu3_mu3_o3
  (
  i0,
  i1,
  o
  );

  input [2:0] i0;
  input [2:0] i1;
  output [2:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_nb0;
  wire net_nb1;
  wire net_nb2;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;

  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b2 (net_nb2, net_b2);

endmodule 

module add_pu4_mu4_o5
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output [4:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_nb0;
  wire net_nb1;
  wire net_nb2;
  wire net_nb3;
  wire net_ncout;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;

  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[4] = net_ncout;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);
  not inv_cout (net_ncout, net_cout3);

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_FADD
  (
  input a,
  input b,
  input c,
  output sum,
  output cout
  );

  wire prop;
  wire not_prop;
  wire sel_i0;
  wire sel_i1;

  xor u0 (prop, a, b);
  xor u1 (sum, prop, c);
  not u2 (not_prop, prop);
  and u3 (sel_i1, prop, c);
  and u4 (sel_i0, not_prop, a);
  or  u5 (cout, sel_i0, sel_i1);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

